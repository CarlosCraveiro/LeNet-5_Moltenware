// parallel.v

// Generated using ACDS version 23.1 991

`timescale 1 ps / 1 ps
module parallel (
		input  wire  clk_clk,                        //                        clk.clk
		input  wire  uart_0_external_connection_rxd, // uart_0_external_connection.rxd
		output wire  uart_0_external_connection_txd  //                           .txd
	);

	wire         hypervisor_debug_reset_request_reset;                                             // hypervisor:debug_reset_request -> rst_controller:reset_in0
	wire         hypervisor_custom_instruction_master_readra;                                      // hypervisor:E_ci_combo_readra -> hypervisor_custom_instruction_master_translator:ci_slave_readra
	wire         hypervisor_custom_instruction_master_readrb;                                      // hypervisor:E_ci_combo_readrb -> hypervisor_custom_instruction_master_translator:ci_slave_readrb
	wire   [4:0] hypervisor_custom_instruction_master_multi_b;                                     // hypervisor:A_ci_multi_b -> hypervisor_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] hypervisor_custom_instruction_master_multi_c;                                     // hypervisor:A_ci_multi_c -> hypervisor_custom_instruction_master_translator:ci_slave_multi_c
	wire         hypervisor_custom_instruction_master_reset_req;                                   // hypervisor:A_ci_multi_reset_req -> hypervisor_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] hypervisor_custom_instruction_master_multi_a;                                     // hypervisor:A_ci_multi_a -> hypervisor_custom_instruction_master_translator:ci_slave_multi_a
	wire  [31:0] hypervisor_custom_instruction_master_result;                                      // hypervisor_custom_instruction_master_translator:ci_slave_result -> hypervisor:E_ci_combo_result
	wire  [31:0] hypervisor_custom_instruction_master_datab;                                       // hypervisor:E_ci_combo_datab -> hypervisor_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] hypervisor_custom_instruction_master_dataa;                                       // hypervisor:E_ci_combo_dataa -> hypervisor_custom_instruction_master_translator:ci_slave_dataa
	wire         hypervisor_custom_instruction_master_writerc;                                     // hypervisor:E_ci_combo_writerc -> hypervisor_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] hypervisor_custom_instruction_master_multi_dataa;                                 // hypervisor:A_ci_multi_dataa -> hypervisor_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         hypervisor_custom_instruction_master_multi_writerc;                               // hypervisor:A_ci_multi_writerc -> hypervisor_custom_instruction_master_translator:ci_slave_multi_writerc
	wire   [4:0] hypervisor_custom_instruction_master_a;                                           // hypervisor:E_ci_combo_a -> hypervisor_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] hypervisor_custom_instruction_master_b;                                           // hypervisor:E_ci_combo_b -> hypervisor_custom_instruction_master_translator:ci_slave_b
	wire  [31:0] hypervisor_custom_instruction_master_multi_result;                                // hypervisor_custom_instruction_master_translator:ci_slave_multi_result -> hypervisor:A_ci_multi_result
	wire         hypervisor_custom_instruction_master_clk;                                         // hypervisor:A_ci_multi_clock -> hypervisor_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] hypervisor_custom_instruction_master_multi_datab;                                 // hypervisor:A_ci_multi_datab -> hypervisor_custom_instruction_master_translator:ci_slave_multi_datab
	wire   [4:0] hypervisor_custom_instruction_master_c;                                           // hypervisor:E_ci_combo_c -> hypervisor_custom_instruction_master_translator:ci_slave_c
	wire  [31:0] hypervisor_custom_instruction_master_ipending;                                    // hypervisor:E_ci_combo_ipending -> hypervisor_custom_instruction_master_translator:ci_slave_ipending
	wire         hypervisor_custom_instruction_master_start;                                       // hypervisor:A_ci_multi_start -> hypervisor_custom_instruction_master_translator:ci_slave_multi_start
	wire         hypervisor_custom_instruction_master_done;                                        // hypervisor_custom_instruction_master_translator:ci_slave_multi_done -> hypervisor:A_ci_multi_done
	wire   [7:0] hypervisor_custom_instruction_master_n;                                           // hypervisor:E_ci_combo_n -> hypervisor_custom_instruction_master_translator:ci_slave_n
	wire         hypervisor_custom_instruction_master_estatus;                                     // hypervisor:E_ci_combo_estatus -> hypervisor_custom_instruction_master_translator:ci_slave_estatus
	wire         hypervisor_custom_instruction_master_clk_en;                                      // hypervisor:A_ci_multi_clk_en -> hypervisor_custom_instruction_master_translator:ci_slave_multi_clken
	wire         hypervisor_custom_instruction_master_reset;                                       // hypervisor:A_ci_multi_reset -> hypervisor_custom_instruction_master_translator:ci_slave_multi_reset
	wire         hypervisor_custom_instruction_master_multi_readrb;                                // hypervisor:A_ci_multi_readrb -> hypervisor_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         hypervisor_custom_instruction_master_multi_readra;                                // hypervisor:A_ci_multi_readra -> hypervisor_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] hypervisor_custom_instruction_master_multi_n;                                     // hypervisor:A_ci_multi_n -> hypervisor_custom_instruction_master_translator:ci_slave_multi_n
	wire  [31:0] hypervisor_custom_instruction_master_translator_comb_ci_master_result;            // hypervisor_custom_instruction_master_comb_xconnect:ci_slave_result -> hypervisor_custom_instruction_master_translator:comb_ci_master_result
	wire         hypervisor_custom_instruction_master_translator_comb_ci_master_readra;            // hypervisor_custom_instruction_master_translator:comb_ci_master_readra -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] hypervisor_custom_instruction_master_translator_comb_ci_master_a;                 // hypervisor_custom_instruction_master_translator:comb_ci_master_a -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] hypervisor_custom_instruction_master_translator_comb_ci_master_b;                 // hypervisor_custom_instruction_master_translator:comb_ci_master_b -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         hypervisor_custom_instruction_master_translator_comb_ci_master_readrb;            // hypervisor_custom_instruction_master_translator:comb_ci_master_readrb -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] hypervisor_custom_instruction_master_translator_comb_ci_master_c;                 // hypervisor_custom_instruction_master_translator:comb_ci_master_c -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         hypervisor_custom_instruction_master_translator_comb_ci_master_estatus;           // hypervisor_custom_instruction_master_translator:comb_ci_master_estatus -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] hypervisor_custom_instruction_master_translator_comb_ci_master_ipending;          // hypervisor_custom_instruction_master_translator:comb_ci_master_ipending -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] hypervisor_custom_instruction_master_translator_comb_ci_master_datab;             // hypervisor_custom_instruction_master_translator:comb_ci_master_datab -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] hypervisor_custom_instruction_master_translator_comb_ci_master_dataa;             // hypervisor_custom_instruction_master_translator:comb_ci_master_dataa -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         hypervisor_custom_instruction_master_translator_comb_ci_master_writerc;           // hypervisor_custom_instruction_master_translator:comb_ci_master_writerc -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] hypervisor_custom_instruction_master_translator_comb_ci_master_n;                 // hypervisor_custom_instruction_master_translator:comb_ci_master_n -> hypervisor_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] hypervisor_custom_instruction_master_comb_xconnect_ci_master0_result;             // hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_result -> hypervisor_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         hypervisor_custom_instruction_master_comb_xconnect_ci_master0_readra;             // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_readra -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] hypervisor_custom_instruction_master_comb_xconnect_ci_master0_a;                  // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_a -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] hypervisor_custom_instruction_master_comb_xconnect_ci_master0_b;                  // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_b -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         hypervisor_custom_instruction_master_comb_xconnect_ci_master0_readrb;             // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_readrb -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] hypervisor_custom_instruction_master_comb_xconnect_ci_master0_c;                  // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_c -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         hypervisor_custom_instruction_master_comb_xconnect_ci_master0_estatus;            // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_estatus -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] hypervisor_custom_instruction_master_comb_xconnect_ci_master0_ipending;           // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_ipending -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] hypervisor_custom_instruction_master_comb_xconnect_ci_master0_datab;              // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_datab -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] hypervisor_custom_instruction_master_comb_xconnect_ci_master0_dataa;              // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_dataa -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         hypervisor_custom_instruction_master_comb_xconnect_ci_master0_writerc;            // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_writerc -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] hypervisor_custom_instruction_master_comb_xconnect_ci_master0_n;                  // hypervisor_custom_instruction_master_comb_xconnect:ci_master0_n -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_result;     // nios2_fpu:s1_result -> hypervisor_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_datab;      // hypervisor_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios2_fpu:s1_datab
	wire  [31:0] hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_dataa;      // hypervisor_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios2_fpu:s1_dataa
	wire   [3:0] hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_n;          // hypervisor_custom_instruction_master_comb_slave_translator0:ci_master_n -> nios2_fpu:s1_n
	wire         hypervisor_custom_instruction_master_translator_multi_ci_master_readra;           // hypervisor_custom_instruction_master_translator:multi_ci_master_readra -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] hypervisor_custom_instruction_master_translator_multi_ci_master_a;                // hypervisor_custom_instruction_master_translator:multi_ci_master_a -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] hypervisor_custom_instruction_master_translator_multi_ci_master_b;                // hypervisor_custom_instruction_master_translator:multi_ci_master_b -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         hypervisor_custom_instruction_master_translator_multi_ci_master_clk;              // hypervisor_custom_instruction_master_translator:multi_ci_master_clk -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         hypervisor_custom_instruction_master_translator_multi_ci_master_readrb;           // hypervisor_custom_instruction_master_translator:multi_ci_master_readrb -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] hypervisor_custom_instruction_master_translator_multi_ci_master_c;                // hypervisor_custom_instruction_master_translator:multi_ci_master_c -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         hypervisor_custom_instruction_master_translator_multi_ci_master_start;            // hypervisor_custom_instruction_master_translator:multi_ci_master_start -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         hypervisor_custom_instruction_master_translator_multi_ci_master_reset_req;        // hypervisor_custom_instruction_master_translator:multi_ci_master_reset_req -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         hypervisor_custom_instruction_master_translator_multi_ci_master_done;             // hypervisor_custom_instruction_master_multi_xconnect:ci_slave_done -> hypervisor_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] hypervisor_custom_instruction_master_translator_multi_ci_master_n;                // hypervisor_custom_instruction_master_translator:multi_ci_master_n -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] hypervisor_custom_instruction_master_translator_multi_ci_master_result;           // hypervisor_custom_instruction_master_multi_xconnect:ci_slave_result -> hypervisor_custom_instruction_master_translator:multi_ci_master_result
	wire         hypervisor_custom_instruction_master_translator_multi_ci_master_clk_en;           // hypervisor_custom_instruction_master_translator:multi_ci_master_clken -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] hypervisor_custom_instruction_master_translator_multi_ci_master_datab;            // hypervisor_custom_instruction_master_translator:multi_ci_master_datab -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] hypervisor_custom_instruction_master_translator_multi_ci_master_dataa;            // hypervisor_custom_instruction_master_translator:multi_ci_master_dataa -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         hypervisor_custom_instruction_master_translator_multi_ci_master_reset;            // hypervisor_custom_instruction_master_translator:multi_ci_master_reset -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         hypervisor_custom_instruction_master_translator_multi_ci_master_writerc;          // hypervisor_custom_instruction_master_translator:multi_ci_master_writerc -> hypervisor_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         hypervisor_custom_instruction_master_multi_xconnect_ci_master0_readra;            // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_readra -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] hypervisor_custom_instruction_master_multi_xconnect_ci_master0_a;                 // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_a -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] hypervisor_custom_instruction_master_multi_xconnect_ci_master0_b;                 // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_b -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         hypervisor_custom_instruction_master_multi_xconnect_ci_master0_readrb;            // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_readrb -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] hypervisor_custom_instruction_master_multi_xconnect_ci_master0_c;                 // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_c -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         hypervisor_custom_instruction_master_multi_xconnect_ci_master0_clk;               // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_clk -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] hypervisor_custom_instruction_master_multi_xconnect_ci_master0_ipending;          // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_ipending -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         hypervisor_custom_instruction_master_multi_xconnect_ci_master0_start;             // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_start -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         hypervisor_custom_instruction_master_multi_xconnect_ci_master0_reset_req;         // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         hypervisor_custom_instruction_master_multi_xconnect_ci_master0_done;              // hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_done -> hypervisor_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] hypervisor_custom_instruction_master_multi_xconnect_ci_master0_n;                 // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_n -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] hypervisor_custom_instruction_master_multi_xconnect_ci_master0_result;            // hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_result -> hypervisor_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         hypervisor_custom_instruction_master_multi_xconnect_ci_master0_estatus;           // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_estatus -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         hypervisor_custom_instruction_master_multi_xconnect_ci_master0_clk_en;            // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_clken -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] hypervisor_custom_instruction_master_multi_xconnect_ci_master0_datab;             // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_datab -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] hypervisor_custom_instruction_master_multi_xconnect_ci_master0_dataa;             // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_dataa -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         hypervisor_custom_instruction_master_multi_xconnect_ci_master0_reset;             // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_reset -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         hypervisor_custom_instruction_master_multi_xconnect_ci_master0_writerc;           // hypervisor_custom_instruction_master_multi_xconnect:ci_master0_writerc -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_result;    // nios2_fpu:s2_result -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_clk;       // hypervisor_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios2_fpu:s2_clk
	wire         hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;    // hypervisor_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios2_fpu:s2_clk_en
	wire  [31:0] hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_datab;     // hypervisor_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios2_fpu:s2_datab
	wire  [31:0] hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_dataa;     // hypervisor_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios2_fpu:s2_dataa
	wire         hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_start;     // hypervisor_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios2_fpu:s2_start
	wire         hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_reset;     // hypervisor_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios2_fpu:s2_reset
	wire         hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_reset_req; // hypervisor_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> nios2_fpu:s2_reset_req
	wire         hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_done;      // nios2_fpu:s2_done -> hypervisor_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_n;         // hypervisor_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios2_fpu:s2_n
	wire         cpu_2_custom_instruction_master_readra;                                           // cpu_2:E_ci_combo_readra -> cpu_2_custom_instruction_master_translator:ci_slave_readra
	wire         cpu_2_custom_instruction_master_readrb;                                           // cpu_2:E_ci_combo_readrb -> cpu_2_custom_instruction_master_translator:ci_slave_readrb
	wire   [4:0] cpu_2_custom_instruction_master_multi_b;                                          // cpu_2:A_ci_multi_b -> cpu_2_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] cpu_2_custom_instruction_master_multi_c;                                          // cpu_2:A_ci_multi_c -> cpu_2_custom_instruction_master_translator:ci_slave_multi_c
	wire         cpu_2_custom_instruction_master_reset_req;                                        // cpu_2:A_ci_multi_reset_req -> cpu_2_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] cpu_2_custom_instruction_master_multi_a;                                          // cpu_2:A_ci_multi_a -> cpu_2_custom_instruction_master_translator:ci_slave_multi_a
	wire  [31:0] cpu_2_custom_instruction_master_result;                                           // cpu_2_custom_instruction_master_translator:ci_slave_result -> cpu_2:E_ci_combo_result
	wire  [31:0] cpu_2_custom_instruction_master_datab;                                            // cpu_2:E_ci_combo_datab -> cpu_2_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] cpu_2_custom_instruction_master_dataa;                                            // cpu_2:E_ci_combo_dataa -> cpu_2_custom_instruction_master_translator:ci_slave_dataa
	wire         cpu_2_custom_instruction_master_writerc;                                          // cpu_2:E_ci_combo_writerc -> cpu_2_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] cpu_2_custom_instruction_master_multi_dataa;                                      // cpu_2:A_ci_multi_dataa -> cpu_2_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         cpu_2_custom_instruction_master_multi_writerc;                                    // cpu_2:A_ci_multi_writerc -> cpu_2_custom_instruction_master_translator:ci_slave_multi_writerc
	wire   [4:0] cpu_2_custom_instruction_master_a;                                                // cpu_2:E_ci_combo_a -> cpu_2_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] cpu_2_custom_instruction_master_b;                                                // cpu_2:E_ci_combo_b -> cpu_2_custom_instruction_master_translator:ci_slave_b
	wire  [31:0] cpu_2_custom_instruction_master_multi_result;                                     // cpu_2_custom_instruction_master_translator:ci_slave_multi_result -> cpu_2:A_ci_multi_result
	wire         cpu_2_custom_instruction_master_clk;                                              // cpu_2:A_ci_multi_clock -> cpu_2_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] cpu_2_custom_instruction_master_multi_datab;                                      // cpu_2:A_ci_multi_datab -> cpu_2_custom_instruction_master_translator:ci_slave_multi_datab
	wire   [4:0] cpu_2_custom_instruction_master_c;                                                // cpu_2:E_ci_combo_c -> cpu_2_custom_instruction_master_translator:ci_slave_c
	wire  [31:0] cpu_2_custom_instruction_master_ipending;                                         // cpu_2:E_ci_combo_ipending -> cpu_2_custom_instruction_master_translator:ci_slave_ipending
	wire         cpu_2_custom_instruction_master_start;                                            // cpu_2:A_ci_multi_start -> cpu_2_custom_instruction_master_translator:ci_slave_multi_start
	wire         cpu_2_custom_instruction_master_done;                                             // cpu_2_custom_instruction_master_translator:ci_slave_multi_done -> cpu_2:A_ci_multi_done
	wire   [7:0] cpu_2_custom_instruction_master_n;                                                // cpu_2:E_ci_combo_n -> cpu_2_custom_instruction_master_translator:ci_slave_n
	wire         cpu_2_custom_instruction_master_estatus;                                          // cpu_2:E_ci_combo_estatus -> cpu_2_custom_instruction_master_translator:ci_slave_estatus
	wire         cpu_2_custom_instruction_master_clk_en;                                           // cpu_2:A_ci_multi_clk_en -> cpu_2_custom_instruction_master_translator:ci_slave_multi_clken
	wire         cpu_2_custom_instruction_master_reset;                                            // cpu_2:A_ci_multi_reset -> cpu_2_custom_instruction_master_translator:ci_slave_multi_reset
	wire         cpu_2_custom_instruction_master_multi_readrb;                                     // cpu_2:A_ci_multi_readrb -> cpu_2_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         cpu_2_custom_instruction_master_multi_readra;                                     // cpu_2:A_ci_multi_readra -> cpu_2_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] cpu_2_custom_instruction_master_multi_n;                                          // cpu_2:A_ci_multi_n -> cpu_2_custom_instruction_master_translator:ci_slave_multi_n
	wire  [31:0] cpu_2_custom_instruction_master_translator_comb_ci_master_result;                 // cpu_2_custom_instruction_master_comb_xconnect:ci_slave_result -> cpu_2_custom_instruction_master_translator:comb_ci_master_result
	wire         cpu_2_custom_instruction_master_translator_comb_ci_master_readra;                 // cpu_2_custom_instruction_master_translator:comb_ci_master_readra -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] cpu_2_custom_instruction_master_translator_comb_ci_master_a;                      // cpu_2_custom_instruction_master_translator:comb_ci_master_a -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] cpu_2_custom_instruction_master_translator_comb_ci_master_b;                      // cpu_2_custom_instruction_master_translator:comb_ci_master_b -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         cpu_2_custom_instruction_master_translator_comb_ci_master_readrb;                 // cpu_2_custom_instruction_master_translator:comb_ci_master_readrb -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] cpu_2_custom_instruction_master_translator_comb_ci_master_c;                      // cpu_2_custom_instruction_master_translator:comb_ci_master_c -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         cpu_2_custom_instruction_master_translator_comb_ci_master_estatus;                // cpu_2_custom_instruction_master_translator:comb_ci_master_estatus -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] cpu_2_custom_instruction_master_translator_comb_ci_master_ipending;               // cpu_2_custom_instruction_master_translator:comb_ci_master_ipending -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] cpu_2_custom_instruction_master_translator_comb_ci_master_datab;                  // cpu_2_custom_instruction_master_translator:comb_ci_master_datab -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] cpu_2_custom_instruction_master_translator_comb_ci_master_dataa;                  // cpu_2_custom_instruction_master_translator:comb_ci_master_dataa -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         cpu_2_custom_instruction_master_translator_comb_ci_master_writerc;                // cpu_2_custom_instruction_master_translator:comb_ci_master_writerc -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] cpu_2_custom_instruction_master_translator_comb_ci_master_n;                      // cpu_2_custom_instruction_master_translator:comb_ci_master_n -> cpu_2_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] cpu_2_custom_instruction_master_comb_xconnect_ci_master0_result;                  // cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_result -> cpu_2_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         cpu_2_custom_instruction_master_comb_xconnect_ci_master0_readra;                  // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_readra -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] cpu_2_custom_instruction_master_comb_xconnect_ci_master0_a;                       // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_a -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] cpu_2_custom_instruction_master_comb_xconnect_ci_master0_b;                       // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_b -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         cpu_2_custom_instruction_master_comb_xconnect_ci_master0_readrb;                  // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_readrb -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] cpu_2_custom_instruction_master_comb_xconnect_ci_master0_c;                       // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_c -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         cpu_2_custom_instruction_master_comb_xconnect_ci_master0_estatus;                 // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_estatus -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] cpu_2_custom_instruction_master_comb_xconnect_ci_master0_ipending;                // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_ipending -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] cpu_2_custom_instruction_master_comb_xconnect_ci_master0_datab;                   // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_datab -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] cpu_2_custom_instruction_master_comb_xconnect_ci_master0_dataa;                   // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_dataa -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         cpu_2_custom_instruction_master_comb_xconnect_ci_master0_writerc;                 // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_writerc -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] cpu_2_custom_instruction_master_comb_xconnect_ci_master0_n;                       // cpu_2_custom_instruction_master_comb_xconnect:ci_master0_n -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_result;          // fpu_2:s1_result -> cpu_2_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_datab;           // cpu_2_custom_instruction_master_comb_slave_translator0:ci_master_datab -> fpu_2:s1_datab
	wire  [31:0] cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_dataa;           // cpu_2_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> fpu_2:s1_dataa
	wire   [3:0] cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_n;               // cpu_2_custom_instruction_master_comb_slave_translator0:ci_master_n -> fpu_2:s1_n
	wire         cpu_2_custom_instruction_master_translator_multi_ci_master_readra;                // cpu_2_custom_instruction_master_translator:multi_ci_master_readra -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] cpu_2_custom_instruction_master_translator_multi_ci_master_a;                     // cpu_2_custom_instruction_master_translator:multi_ci_master_a -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] cpu_2_custom_instruction_master_translator_multi_ci_master_b;                     // cpu_2_custom_instruction_master_translator:multi_ci_master_b -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         cpu_2_custom_instruction_master_translator_multi_ci_master_clk;                   // cpu_2_custom_instruction_master_translator:multi_ci_master_clk -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         cpu_2_custom_instruction_master_translator_multi_ci_master_readrb;                // cpu_2_custom_instruction_master_translator:multi_ci_master_readrb -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] cpu_2_custom_instruction_master_translator_multi_ci_master_c;                     // cpu_2_custom_instruction_master_translator:multi_ci_master_c -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         cpu_2_custom_instruction_master_translator_multi_ci_master_start;                 // cpu_2_custom_instruction_master_translator:multi_ci_master_start -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         cpu_2_custom_instruction_master_translator_multi_ci_master_reset_req;             // cpu_2_custom_instruction_master_translator:multi_ci_master_reset_req -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         cpu_2_custom_instruction_master_translator_multi_ci_master_done;                  // cpu_2_custom_instruction_master_multi_xconnect:ci_slave_done -> cpu_2_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] cpu_2_custom_instruction_master_translator_multi_ci_master_n;                     // cpu_2_custom_instruction_master_translator:multi_ci_master_n -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] cpu_2_custom_instruction_master_translator_multi_ci_master_result;                // cpu_2_custom_instruction_master_multi_xconnect:ci_slave_result -> cpu_2_custom_instruction_master_translator:multi_ci_master_result
	wire         cpu_2_custom_instruction_master_translator_multi_ci_master_clk_en;                // cpu_2_custom_instruction_master_translator:multi_ci_master_clken -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] cpu_2_custom_instruction_master_translator_multi_ci_master_datab;                 // cpu_2_custom_instruction_master_translator:multi_ci_master_datab -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] cpu_2_custom_instruction_master_translator_multi_ci_master_dataa;                 // cpu_2_custom_instruction_master_translator:multi_ci_master_dataa -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         cpu_2_custom_instruction_master_translator_multi_ci_master_reset;                 // cpu_2_custom_instruction_master_translator:multi_ci_master_reset -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         cpu_2_custom_instruction_master_translator_multi_ci_master_writerc;               // cpu_2_custom_instruction_master_translator:multi_ci_master_writerc -> cpu_2_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         cpu_2_custom_instruction_master_multi_xconnect_ci_master0_readra;                 // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_readra -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] cpu_2_custom_instruction_master_multi_xconnect_ci_master0_a;                      // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_a -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] cpu_2_custom_instruction_master_multi_xconnect_ci_master0_b;                      // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_b -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         cpu_2_custom_instruction_master_multi_xconnect_ci_master0_readrb;                 // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_readrb -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] cpu_2_custom_instruction_master_multi_xconnect_ci_master0_c;                      // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_c -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         cpu_2_custom_instruction_master_multi_xconnect_ci_master0_clk;                    // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_clk -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] cpu_2_custom_instruction_master_multi_xconnect_ci_master0_ipending;               // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_ipending -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         cpu_2_custom_instruction_master_multi_xconnect_ci_master0_start;                  // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_start -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         cpu_2_custom_instruction_master_multi_xconnect_ci_master0_reset_req;              // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         cpu_2_custom_instruction_master_multi_xconnect_ci_master0_done;                   // cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_done -> cpu_2_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] cpu_2_custom_instruction_master_multi_xconnect_ci_master0_n;                      // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_n -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] cpu_2_custom_instruction_master_multi_xconnect_ci_master0_result;                 // cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_result -> cpu_2_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         cpu_2_custom_instruction_master_multi_xconnect_ci_master0_estatus;                // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_estatus -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         cpu_2_custom_instruction_master_multi_xconnect_ci_master0_clk_en;                 // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_clken -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] cpu_2_custom_instruction_master_multi_xconnect_ci_master0_datab;                  // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_datab -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] cpu_2_custom_instruction_master_multi_xconnect_ci_master0_dataa;                  // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_dataa -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         cpu_2_custom_instruction_master_multi_xconnect_ci_master0_reset;                  // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_reset -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         cpu_2_custom_instruction_master_multi_xconnect_ci_master0_writerc;                // cpu_2_custom_instruction_master_multi_xconnect:ci_master0_writerc -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_result;         // fpu_2:s2_result -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_clk;            // cpu_2_custom_instruction_master_multi_slave_translator0:ci_master_clk -> fpu_2:s2_clk
	wire         cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;         // cpu_2_custom_instruction_master_multi_slave_translator0:ci_master_clken -> fpu_2:s2_clk_en
	wire  [31:0] cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_datab;          // cpu_2_custom_instruction_master_multi_slave_translator0:ci_master_datab -> fpu_2:s2_datab
	wire  [31:0] cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_dataa;          // cpu_2_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> fpu_2:s2_dataa
	wire         cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_start;          // cpu_2_custom_instruction_master_multi_slave_translator0:ci_master_start -> fpu_2:s2_start
	wire         cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_reset;          // cpu_2_custom_instruction_master_multi_slave_translator0:ci_master_reset -> fpu_2:s2_reset
	wire         cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_reset_req;      // cpu_2_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> fpu_2:s2_reset_req
	wire         cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_done;           // fpu_2:s2_done -> cpu_2_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_n;              // cpu_2_custom_instruction_master_multi_slave_translator0:ci_master_n -> fpu_2:s2_n
	wire         cpu_3_custom_instruction_master_readra;                                           // cpu_3:E_ci_combo_readra -> cpu_3_custom_instruction_master_translator:ci_slave_readra
	wire         cpu_3_custom_instruction_master_readrb;                                           // cpu_3:E_ci_combo_readrb -> cpu_3_custom_instruction_master_translator:ci_slave_readrb
	wire   [4:0] cpu_3_custom_instruction_master_multi_b;                                          // cpu_3:A_ci_multi_b -> cpu_3_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] cpu_3_custom_instruction_master_multi_c;                                          // cpu_3:A_ci_multi_c -> cpu_3_custom_instruction_master_translator:ci_slave_multi_c
	wire         cpu_3_custom_instruction_master_reset_req;                                        // cpu_3:A_ci_multi_reset_req -> cpu_3_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] cpu_3_custom_instruction_master_multi_a;                                          // cpu_3:A_ci_multi_a -> cpu_3_custom_instruction_master_translator:ci_slave_multi_a
	wire  [31:0] cpu_3_custom_instruction_master_result;                                           // cpu_3_custom_instruction_master_translator:ci_slave_result -> cpu_3:E_ci_combo_result
	wire  [31:0] cpu_3_custom_instruction_master_datab;                                            // cpu_3:E_ci_combo_datab -> cpu_3_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] cpu_3_custom_instruction_master_dataa;                                            // cpu_3:E_ci_combo_dataa -> cpu_3_custom_instruction_master_translator:ci_slave_dataa
	wire         cpu_3_custom_instruction_master_writerc;                                          // cpu_3:E_ci_combo_writerc -> cpu_3_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] cpu_3_custom_instruction_master_multi_dataa;                                      // cpu_3:A_ci_multi_dataa -> cpu_3_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         cpu_3_custom_instruction_master_multi_writerc;                                    // cpu_3:A_ci_multi_writerc -> cpu_3_custom_instruction_master_translator:ci_slave_multi_writerc
	wire   [4:0] cpu_3_custom_instruction_master_a;                                                // cpu_3:E_ci_combo_a -> cpu_3_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] cpu_3_custom_instruction_master_b;                                                // cpu_3:E_ci_combo_b -> cpu_3_custom_instruction_master_translator:ci_slave_b
	wire  [31:0] cpu_3_custom_instruction_master_multi_result;                                     // cpu_3_custom_instruction_master_translator:ci_slave_multi_result -> cpu_3:A_ci_multi_result
	wire         cpu_3_custom_instruction_master_clk;                                              // cpu_3:A_ci_multi_clock -> cpu_3_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] cpu_3_custom_instruction_master_multi_datab;                                      // cpu_3:A_ci_multi_datab -> cpu_3_custom_instruction_master_translator:ci_slave_multi_datab
	wire   [4:0] cpu_3_custom_instruction_master_c;                                                // cpu_3:E_ci_combo_c -> cpu_3_custom_instruction_master_translator:ci_slave_c
	wire  [31:0] cpu_3_custom_instruction_master_ipending;                                         // cpu_3:E_ci_combo_ipending -> cpu_3_custom_instruction_master_translator:ci_slave_ipending
	wire         cpu_3_custom_instruction_master_start;                                            // cpu_3:A_ci_multi_start -> cpu_3_custom_instruction_master_translator:ci_slave_multi_start
	wire         cpu_3_custom_instruction_master_done;                                             // cpu_3_custom_instruction_master_translator:ci_slave_multi_done -> cpu_3:A_ci_multi_done
	wire   [7:0] cpu_3_custom_instruction_master_n;                                                // cpu_3:E_ci_combo_n -> cpu_3_custom_instruction_master_translator:ci_slave_n
	wire         cpu_3_custom_instruction_master_estatus;                                          // cpu_3:E_ci_combo_estatus -> cpu_3_custom_instruction_master_translator:ci_slave_estatus
	wire         cpu_3_custom_instruction_master_clk_en;                                           // cpu_3:A_ci_multi_clk_en -> cpu_3_custom_instruction_master_translator:ci_slave_multi_clken
	wire         cpu_3_custom_instruction_master_reset;                                            // cpu_3:A_ci_multi_reset -> cpu_3_custom_instruction_master_translator:ci_slave_multi_reset
	wire         cpu_3_custom_instruction_master_multi_readrb;                                     // cpu_3:A_ci_multi_readrb -> cpu_3_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         cpu_3_custom_instruction_master_multi_readra;                                     // cpu_3:A_ci_multi_readra -> cpu_3_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] cpu_3_custom_instruction_master_multi_n;                                          // cpu_3:A_ci_multi_n -> cpu_3_custom_instruction_master_translator:ci_slave_multi_n
	wire  [31:0] cpu_3_custom_instruction_master_translator_comb_ci_master_result;                 // cpu_3_custom_instruction_master_comb_xconnect:ci_slave_result -> cpu_3_custom_instruction_master_translator:comb_ci_master_result
	wire         cpu_3_custom_instruction_master_translator_comb_ci_master_readra;                 // cpu_3_custom_instruction_master_translator:comb_ci_master_readra -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] cpu_3_custom_instruction_master_translator_comb_ci_master_a;                      // cpu_3_custom_instruction_master_translator:comb_ci_master_a -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] cpu_3_custom_instruction_master_translator_comb_ci_master_b;                      // cpu_3_custom_instruction_master_translator:comb_ci_master_b -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         cpu_3_custom_instruction_master_translator_comb_ci_master_readrb;                 // cpu_3_custom_instruction_master_translator:comb_ci_master_readrb -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] cpu_3_custom_instruction_master_translator_comb_ci_master_c;                      // cpu_3_custom_instruction_master_translator:comb_ci_master_c -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         cpu_3_custom_instruction_master_translator_comb_ci_master_estatus;                // cpu_3_custom_instruction_master_translator:comb_ci_master_estatus -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] cpu_3_custom_instruction_master_translator_comb_ci_master_ipending;               // cpu_3_custom_instruction_master_translator:comb_ci_master_ipending -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] cpu_3_custom_instruction_master_translator_comb_ci_master_datab;                  // cpu_3_custom_instruction_master_translator:comb_ci_master_datab -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] cpu_3_custom_instruction_master_translator_comb_ci_master_dataa;                  // cpu_3_custom_instruction_master_translator:comb_ci_master_dataa -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         cpu_3_custom_instruction_master_translator_comb_ci_master_writerc;                // cpu_3_custom_instruction_master_translator:comb_ci_master_writerc -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] cpu_3_custom_instruction_master_translator_comb_ci_master_n;                      // cpu_3_custom_instruction_master_translator:comb_ci_master_n -> cpu_3_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] cpu_3_custom_instruction_master_comb_xconnect_ci_master0_result;                  // cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_result -> cpu_3_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         cpu_3_custom_instruction_master_comb_xconnect_ci_master0_readra;                  // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_readra -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] cpu_3_custom_instruction_master_comb_xconnect_ci_master0_a;                       // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_a -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] cpu_3_custom_instruction_master_comb_xconnect_ci_master0_b;                       // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_b -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         cpu_3_custom_instruction_master_comb_xconnect_ci_master0_readrb;                  // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_readrb -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] cpu_3_custom_instruction_master_comb_xconnect_ci_master0_c;                       // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_c -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         cpu_3_custom_instruction_master_comb_xconnect_ci_master0_estatus;                 // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_estatus -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] cpu_3_custom_instruction_master_comb_xconnect_ci_master0_ipending;                // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_ipending -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] cpu_3_custom_instruction_master_comb_xconnect_ci_master0_datab;                   // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_datab -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] cpu_3_custom_instruction_master_comb_xconnect_ci_master0_dataa;                   // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_dataa -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         cpu_3_custom_instruction_master_comb_xconnect_ci_master0_writerc;                 // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_writerc -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] cpu_3_custom_instruction_master_comb_xconnect_ci_master0_n;                       // cpu_3_custom_instruction_master_comb_xconnect:ci_master0_n -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_result;          // fpu_3:s1_result -> cpu_3_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_datab;           // cpu_3_custom_instruction_master_comb_slave_translator0:ci_master_datab -> fpu_3:s1_datab
	wire  [31:0] cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_dataa;           // cpu_3_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> fpu_3:s1_dataa
	wire   [3:0] cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_n;               // cpu_3_custom_instruction_master_comb_slave_translator0:ci_master_n -> fpu_3:s1_n
	wire         cpu_3_custom_instruction_master_translator_multi_ci_master_readra;                // cpu_3_custom_instruction_master_translator:multi_ci_master_readra -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] cpu_3_custom_instruction_master_translator_multi_ci_master_a;                     // cpu_3_custom_instruction_master_translator:multi_ci_master_a -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] cpu_3_custom_instruction_master_translator_multi_ci_master_b;                     // cpu_3_custom_instruction_master_translator:multi_ci_master_b -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         cpu_3_custom_instruction_master_translator_multi_ci_master_clk;                   // cpu_3_custom_instruction_master_translator:multi_ci_master_clk -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         cpu_3_custom_instruction_master_translator_multi_ci_master_readrb;                // cpu_3_custom_instruction_master_translator:multi_ci_master_readrb -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] cpu_3_custom_instruction_master_translator_multi_ci_master_c;                     // cpu_3_custom_instruction_master_translator:multi_ci_master_c -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         cpu_3_custom_instruction_master_translator_multi_ci_master_start;                 // cpu_3_custom_instruction_master_translator:multi_ci_master_start -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         cpu_3_custom_instruction_master_translator_multi_ci_master_reset_req;             // cpu_3_custom_instruction_master_translator:multi_ci_master_reset_req -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         cpu_3_custom_instruction_master_translator_multi_ci_master_done;                  // cpu_3_custom_instruction_master_multi_xconnect:ci_slave_done -> cpu_3_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] cpu_3_custom_instruction_master_translator_multi_ci_master_n;                     // cpu_3_custom_instruction_master_translator:multi_ci_master_n -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] cpu_3_custom_instruction_master_translator_multi_ci_master_result;                // cpu_3_custom_instruction_master_multi_xconnect:ci_slave_result -> cpu_3_custom_instruction_master_translator:multi_ci_master_result
	wire         cpu_3_custom_instruction_master_translator_multi_ci_master_clk_en;                // cpu_3_custom_instruction_master_translator:multi_ci_master_clken -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] cpu_3_custom_instruction_master_translator_multi_ci_master_datab;                 // cpu_3_custom_instruction_master_translator:multi_ci_master_datab -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] cpu_3_custom_instruction_master_translator_multi_ci_master_dataa;                 // cpu_3_custom_instruction_master_translator:multi_ci_master_dataa -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         cpu_3_custom_instruction_master_translator_multi_ci_master_reset;                 // cpu_3_custom_instruction_master_translator:multi_ci_master_reset -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         cpu_3_custom_instruction_master_translator_multi_ci_master_writerc;               // cpu_3_custom_instruction_master_translator:multi_ci_master_writerc -> cpu_3_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         cpu_3_custom_instruction_master_multi_xconnect_ci_master0_readra;                 // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_readra -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] cpu_3_custom_instruction_master_multi_xconnect_ci_master0_a;                      // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_a -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] cpu_3_custom_instruction_master_multi_xconnect_ci_master0_b;                      // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_b -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         cpu_3_custom_instruction_master_multi_xconnect_ci_master0_readrb;                 // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_readrb -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] cpu_3_custom_instruction_master_multi_xconnect_ci_master0_c;                      // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_c -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         cpu_3_custom_instruction_master_multi_xconnect_ci_master0_clk;                    // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_clk -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] cpu_3_custom_instruction_master_multi_xconnect_ci_master0_ipending;               // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_ipending -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         cpu_3_custom_instruction_master_multi_xconnect_ci_master0_start;                  // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_start -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         cpu_3_custom_instruction_master_multi_xconnect_ci_master0_reset_req;              // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         cpu_3_custom_instruction_master_multi_xconnect_ci_master0_done;                   // cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_done -> cpu_3_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] cpu_3_custom_instruction_master_multi_xconnect_ci_master0_n;                      // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_n -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] cpu_3_custom_instruction_master_multi_xconnect_ci_master0_result;                 // cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_result -> cpu_3_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         cpu_3_custom_instruction_master_multi_xconnect_ci_master0_estatus;                // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_estatus -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         cpu_3_custom_instruction_master_multi_xconnect_ci_master0_clk_en;                 // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_clken -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] cpu_3_custom_instruction_master_multi_xconnect_ci_master0_datab;                  // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_datab -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] cpu_3_custom_instruction_master_multi_xconnect_ci_master0_dataa;                  // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_dataa -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         cpu_3_custom_instruction_master_multi_xconnect_ci_master0_reset;                  // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_reset -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         cpu_3_custom_instruction_master_multi_xconnect_ci_master0_writerc;                // cpu_3_custom_instruction_master_multi_xconnect:ci_master0_writerc -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_result;         // fpu_3:s2_result -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_clk;            // cpu_3_custom_instruction_master_multi_slave_translator0:ci_master_clk -> fpu_3:s2_clk
	wire         cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;         // cpu_3_custom_instruction_master_multi_slave_translator0:ci_master_clken -> fpu_3:s2_clk_en
	wire  [31:0] cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_datab;          // cpu_3_custom_instruction_master_multi_slave_translator0:ci_master_datab -> fpu_3:s2_datab
	wire  [31:0] cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_dataa;          // cpu_3_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> fpu_3:s2_dataa
	wire         cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_start;          // cpu_3_custom_instruction_master_multi_slave_translator0:ci_master_start -> fpu_3:s2_start
	wire         cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_reset;          // cpu_3_custom_instruction_master_multi_slave_translator0:ci_master_reset -> fpu_3:s2_reset
	wire         cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_reset_req;      // cpu_3_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> fpu_3:s2_reset_req
	wire         cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_done;           // fpu_3:s2_done -> cpu_3_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_n;              // cpu_3_custom_instruction_master_multi_slave_translator0:ci_master_n -> fpu_3:s2_n
	wire         cpu_0_custom_instruction_master_readra;                                           // cpu_0:E_ci_combo_readra -> cpu_0_custom_instruction_master_translator:ci_slave_readra
	wire         cpu_0_custom_instruction_master_readrb;                                           // cpu_0:E_ci_combo_readrb -> cpu_0_custom_instruction_master_translator:ci_slave_readrb
	wire   [4:0] cpu_0_custom_instruction_master_multi_b;                                          // cpu_0:A_ci_multi_b -> cpu_0_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] cpu_0_custom_instruction_master_multi_c;                                          // cpu_0:A_ci_multi_c -> cpu_0_custom_instruction_master_translator:ci_slave_multi_c
	wire         cpu_0_custom_instruction_master_reset_req;                                        // cpu_0:A_ci_multi_reset_req -> cpu_0_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] cpu_0_custom_instruction_master_multi_a;                                          // cpu_0:A_ci_multi_a -> cpu_0_custom_instruction_master_translator:ci_slave_multi_a
	wire  [31:0] cpu_0_custom_instruction_master_result;                                           // cpu_0_custom_instruction_master_translator:ci_slave_result -> cpu_0:E_ci_combo_result
	wire  [31:0] cpu_0_custom_instruction_master_datab;                                            // cpu_0:E_ci_combo_datab -> cpu_0_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] cpu_0_custom_instruction_master_dataa;                                            // cpu_0:E_ci_combo_dataa -> cpu_0_custom_instruction_master_translator:ci_slave_dataa
	wire         cpu_0_custom_instruction_master_writerc;                                          // cpu_0:E_ci_combo_writerc -> cpu_0_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] cpu_0_custom_instruction_master_multi_dataa;                                      // cpu_0:A_ci_multi_dataa -> cpu_0_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         cpu_0_custom_instruction_master_multi_writerc;                                    // cpu_0:A_ci_multi_writerc -> cpu_0_custom_instruction_master_translator:ci_slave_multi_writerc
	wire   [4:0] cpu_0_custom_instruction_master_a;                                                // cpu_0:E_ci_combo_a -> cpu_0_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] cpu_0_custom_instruction_master_b;                                                // cpu_0:E_ci_combo_b -> cpu_0_custom_instruction_master_translator:ci_slave_b
	wire  [31:0] cpu_0_custom_instruction_master_multi_result;                                     // cpu_0_custom_instruction_master_translator:ci_slave_multi_result -> cpu_0:A_ci_multi_result
	wire         cpu_0_custom_instruction_master_clk;                                              // cpu_0:A_ci_multi_clock -> cpu_0_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] cpu_0_custom_instruction_master_multi_datab;                                      // cpu_0:A_ci_multi_datab -> cpu_0_custom_instruction_master_translator:ci_slave_multi_datab
	wire   [4:0] cpu_0_custom_instruction_master_c;                                                // cpu_0:E_ci_combo_c -> cpu_0_custom_instruction_master_translator:ci_slave_c
	wire  [31:0] cpu_0_custom_instruction_master_ipending;                                         // cpu_0:E_ci_combo_ipending -> cpu_0_custom_instruction_master_translator:ci_slave_ipending
	wire         cpu_0_custom_instruction_master_start;                                            // cpu_0:A_ci_multi_start -> cpu_0_custom_instruction_master_translator:ci_slave_multi_start
	wire         cpu_0_custom_instruction_master_done;                                             // cpu_0_custom_instruction_master_translator:ci_slave_multi_done -> cpu_0:A_ci_multi_done
	wire   [7:0] cpu_0_custom_instruction_master_n;                                                // cpu_0:E_ci_combo_n -> cpu_0_custom_instruction_master_translator:ci_slave_n
	wire         cpu_0_custom_instruction_master_estatus;                                          // cpu_0:E_ci_combo_estatus -> cpu_0_custom_instruction_master_translator:ci_slave_estatus
	wire         cpu_0_custom_instruction_master_clk_en;                                           // cpu_0:A_ci_multi_clk_en -> cpu_0_custom_instruction_master_translator:ci_slave_multi_clken
	wire         cpu_0_custom_instruction_master_reset;                                            // cpu_0:A_ci_multi_reset -> cpu_0_custom_instruction_master_translator:ci_slave_multi_reset
	wire         cpu_0_custom_instruction_master_multi_readrb;                                     // cpu_0:A_ci_multi_readrb -> cpu_0_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         cpu_0_custom_instruction_master_multi_readra;                                     // cpu_0:A_ci_multi_readra -> cpu_0_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] cpu_0_custom_instruction_master_multi_n;                                          // cpu_0:A_ci_multi_n -> cpu_0_custom_instruction_master_translator:ci_slave_multi_n
	wire  [31:0] cpu_0_custom_instruction_master_translator_comb_ci_master_result;                 // cpu_0_custom_instruction_master_comb_xconnect:ci_slave_result -> cpu_0_custom_instruction_master_translator:comb_ci_master_result
	wire         cpu_0_custom_instruction_master_translator_comb_ci_master_readra;                 // cpu_0_custom_instruction_master_translator:comb_ci_master_readra -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] cpu_0_custom_instruction_master_translator_comb_ci_master_a;                      // cpu_0_custom_instruction_master_translator:comb_ci_master_a -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] cpu_0_custom_instruction_master_translator_comb_ci_master_b;                      // cpu_0_custom_instruction_master_translator:comb_ci_master_b -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         cpu_0_custom_instruction_master_translator_comb_ci_master_readrb;                 // cpu_0_custom_instruction_master_translator:comb_ci_master_readrb -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] cpu_0_custom_instruction_master_translator_comb_ci_master_c;                      // cpu_0_custom_instruction_master_translator:comb_ci_master_c -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         cpu_0_custom_instruction_master_translator_comb_ci_master_estatus;                // cpu_0_custom_instruction_master_translator:comb_ci_master_estatus -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] cpu_0_custom_instruction_master_translator_comb_ci_master_ipending;               // cpu_0_custom_instruction_master_translator:comb_ci_master_ipending -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] cpu_0_custom_instruction_master_translator_comb_ci_master_datab;                  // cpu_0_custom_instruction_master_translator:comb_ci_master_datab -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] cpu_0_custom_instruction_master_translator_comb_ci_master_dataa;                  // cpu_0_custom_instruction_master_translator:comb_ci_master_dataa -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         cpu_0_custom_instruction_master_translator_comb_ci_master_writerc;                // cpu_0_custom_instruction_master_translator:comb_ci_master_writerc -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] cpu_0_custom_instruction_master_translator_comb_ci_master_n;                      // cpu_0_custom_instruction_master_translator:comb_ci_master_n -> cpu_0_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] cpu_0_custom_instruction_master_comb_xconnect_ci_master0_result;                  // cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_result -> cpu_0_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         cpu_0_custom_instruction_master_comb_xconnect_ci_master0_readra;                  // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_readra -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] cpu_0_custom_instruction_master_comb_xconnect_ci_master0_a;                       // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_a -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] cpu_0_custom_instruction_master_comb_xconnect_ci_master0_b;                       // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_b -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         cpu_0_custom_instruction_master_comb_xconnect_ci_master0_readrb;                  // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_readrb -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] cpu_0_custom_instruction_master_comb_xconnect_ci_master0_c;                       // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_c -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         cpu_0_custom_instruction_master_comb_xconnect_ci_master0_estatus;                 // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_estatus -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] cpu_0_custom_instruction_master_comb_xconnect_ci_master0_ipending;                // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_ipending -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] cpu_0_custom_instruction_master_comb_xconnect_ci_master0_datab;                   // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_datab -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] cpu_0_custom_instruction_master_comb_xconnect_ci_master0_dataa;                   // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_dataa -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         cpu_0_custom_instruction_master_comb_xconnect_ci_master0_writerc;                 // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_writerc -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] cpu_0_custom_instruction_master_comb_xconnect_ci_master0_n;                       // cpu_0_custom_instruction_master_comb_xconnect:ci_master0_n -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_result;          // fpu_0:s1_result -> cpu_0_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_datab;           // cpu_0_custom_instruction_master_comb_slave_translator0:ci_master_datab -> fpu_0:s1_datab
	wire  [31:0] cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa;           // cpu_0_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> fpu_0:s1_dataa
	wire   [3:0] cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_n;               // cpu_0_custom_instruction_master_comb_slave_translator0:ci_master_n -> fpu_0:s1_n
	wire         cpu_0_custom_instruction_master_translator_multi_ci_master_readra;                // cpu_0_custom_instruction_master_translator:multi_ci_master_readra -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] cpu_0_custom_instruction_master_translator_multi_ci_master_a;                     // cpu_0_custom_instruction_master_translator:multi_ci_master_a -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] cpu_0_custom_instruction_master_translator_multi_ci_master_b;                     // cpu_0_custom_instruction_master_translator:multi_ci_master_b -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         cpu_0_custom_instruction_master_translator_multi_ci_master_clk;                   // cpu_0_custom_instruction_master_translator:multi_ci_master_clk -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         cpu_0_custom_instruction_master_translator_multi_ci_master_readrb;                // cpu_0_custom_instruction_master_translator:multi_ci_master_readrb -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] cpu_0_custom_instruction_master_translator_multi_ci_master_c;                     // cpu_0_custom_instruction_master_translator:multi_ci_master_c -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         cpu_0_custom_instruction_master_translator_multi_ci_master_start;                 // cpu_0_custom_instruction_master_translator:multi_ci_master_start -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         cpu_0_custom_instruction_master_translator_multi_ci_master_reset_req;             // cpu_0_custom_instruction_master_translator:multi_ci_master_reset_req -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         cpu_0_custom_instruction_master_translator_multi_ci_master_done;                  // cpu_0_custom_instruction_master_multi_xconnect:ci_slave_done -> cpu_0_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] cpu_0_custom_instruction_master_translator_multi_ci_master_n;                     // cpu_0_custom_instruction_master_translator:multi_ci_master_n -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] cpu_0_custom_instruction_master_translator_multi_ci_master_result;                // cpu_0_custom_instruction_master_multi_xconnect:ci_slave_result -> cpu_0_custom_instruction_master_translator:multi_ci_master_result
	wire         cpu_0_custom_instruction_master_translator_multi_ci_master_clk_en;                // cpu_0_custom_instruction_master_translator:multi_ci_master_clken -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] cpu_0_custom_instruction_master_translator_multi_ci_master_datab;                 // cpu_0_custom_instruction_master_translator:multi_ci_master_datab -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] cpu_0_custom_instruction_master_translator_multi_ci_master_dataa;                 // cpu_0_custom_instruction_master_translator:multi_ci_master_dataa -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         cpu_0_custom_instruction_master_translator_multi_ci_master_reset;                 // cpu_0_custom_instruction_master_translator:multi_ci_master_reset -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         cpu_0_custom_instruction_master_translator_multi_ci_master_writerc;               // cpu_0_custom_instruction_master_translator:multi_ci_master_writerc -> cpu_0_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         cpu_0_custom_instruction_master_multi_xconnect_ci_master0_readra;                 // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_readra -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] cpu_0_custom_instruction_master_multi_xconnect_ci_master0_a;                      // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_a -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] cpu_0_custom_instruction_master_multi_xconnect_ci_master0_b;                      // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_b -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         cpu_0_custom_instruction_master_multi_xconnect_ci_master0_readrb;                 // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_readrb -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] cpu_0_custom_instruction_master_multi_xconnect_ci_master0_c;                      // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_c -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         cpu_0_custom_instruction_master_multi_xconnect_ci_master0_clk;                    // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_clk -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] cpu_0_custom_instruction_master_multi_xconnect_ci_master0_ipending;               // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_ipending -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         cpu_0_custom_instruction_master_multi_xconnect_ci_master0_start;                  // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_start -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         cpu_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req;              // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         cpu_0_custom_instruction_master_multi_xconnect_ci_master0_done;                   // cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_done -> cpu_0_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] cpu_0_custom_instruction_master_multi_xconnect_ci_master0_n;                      // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_n -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] cpu_0_custom_instruction_master_multi_xconnect_ci_master0_result;                 // cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_result -> cpu_0_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         cpu_0_custom_instruction_master_multi_xconnect_ci_master0_estatus;                // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_estatus -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         cpu_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en;                 // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_clken -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] cpu_0_custom_instruction_master_multi_xconnect_ci_master0_datab;                  // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_datab -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] cpu_0_custom_instruction_master_multi_xconnect_ci_master0_dataa;                  // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_dataa -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         cpu_0_custom_instruction_master_multi_xconnect_ci_master0_reset;                  // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_reset -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         cpu_0_custom_instruction_master_multi_xconnect_ci_master0_writerc;                // cpu_0_custom_instruction_master_multi_xconnect:ci_master0_writerc -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_result;         // fpu_0:s2_result -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_clk;            // cpu_0_custom_instruction_master_multi_slave_translator0:ci_master_clk -> fpu_0:s2_clk
	wire         cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;         // cpu_0_custom_instruction_master_multi_slave_translator0:ci_master_clken -> fpu_0:s2_clk_en
	wire  [31:0] cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_datab;          // cpu_0_custom_instruction_master_multi_slave_translator0:ci_master_datab -> fpu_0:s2_datab
	wire  [31:0] cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa;          // cpu_0_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> fpu_0:s2_dataa
	wire         cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_start;          // cpu_0_custom_instruction_master_multi_slave_translator0:ci_master_start -> fpu_0:s2_start
	wire         cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_reset;          // cpu_0_custom_instruction_master_multi_slave_translator0:ci_master_reset -> fpu_0:s2_reset
	wire         cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_reset_req;      // cpu_0_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> fpu_0:s2_reset_req
	wire         cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_done;           // fpu_0:s2_done -> cpu_0_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_n;              // cpu_0_custom_instruction_master_multi_slave_translator0:ci_master_n -> fpu_0:s2_n
	wire  [31:0] hypervisor_data_master_readdata;                                                  // mm_interconnect_0:hypervisor_data_master_readdata -> hypervisor:d_readdata
	wire         hypervisor_data_master_waitrequest;                                               // mm_interconnect_0:hypervisor_data_master_waitrequest -> hypervisor:d_waitrequest
	wire         hypervisor_data_master_debugaccess;                                               // hypervisor:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:hypervisor_data_master_debugaccess
	wire  [22:0] hypervisor_data_master_address;                                                   // hypervisor:d_address -> mm_interconnect_0:hypervisor_data_master_address
	wire   [3:0] hypervisor_data_master_byteenable;                                                // hypervisor:d_byteenable -> mm_interconnect_0:hypervisor_data_master_byteenable
	wire         hypervisor_data_master_read;                                                      // hypervisor:d_read -> mm_interconnect_0:hypervisor_data_master_read
	wire         hypervisor_data_master_readdatavalid;                                             // mm_interconnect_0:hypervisor_data_master_readdatavalid -> hypervisor:d_readdatavalid
	wire         hypervisor_data_master_write;                                                     // hypervisor:d_write -> mm_interconnect_0:hypervisor_data_master_write
	wire  [31:0] hypervisor_data_master_writedata;                                                 // hypervisor:d_writedata -> mm_interconnect_0:hypervisor_data_master_writedata
	wire  [31:0] cpu_0_data_master_readdata;                                                       // mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_waitrequest;                                                    // mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	wire         cpu_0_data_master_debugaccess;                                                    // cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	wire  [22:0] cpu_0_data_master_address;                                                        // cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	wire   [3:0] cpu_0_data_master_byteenable;                                                     // cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	wire         cpu_0_data_master_read;                                                           // cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	wire         cpu_0_data_master_readdatavalid;                                                  // mm_interconnect_0:cpu_0_data_master_readdatavalid -> cpu_0:d_readdatavalid
	wire         cpu_0_data_master_write;                                                          // cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	wire  [31:0] cpu_0_data_master_writedata;                                                      // cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	wire  [31:0] hypervisor_instruction_master_readdata;                                           // mm_interconnect_0:hypervisor_instruction_master_readdata -> hypervisor:i_readdata
	wire         hypervisor_instruction_master_waitrequest;                                        // mm_interconnect_0:hypervisor_instruction_master_waitrequest -> hypervisor:i_waitrequest
	wire  [22:0] hypervisor_instruction_master_address;                                            // hypervisor:i_address -> mm_interconnect_0:hypervisor_instruction_master_address
	wire         hypervisor_instruction_master_read;                                               // hypervisor:i_read -> mm_interconnect_0:hypervisor_instruction_master_read
	wire         hypervisor_instruction_master_readdatavalid;                                      // mm_interconnect_0:hypervisor_instruction_master_readdatavalid -> hypervisor:i_readdatavalid
	wire  [31:0] cpu_0_instruction_master_readdata;                                                // mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	wire         cpu_0_instruction_master_waitrequest;                                             // mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	wire  [22:0] cpu_0_instruction_master_address;                                                 // cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	wire         cpu_0_instruction_master_read;                                                    // cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	wire         cpu_0_instruction_master_readdatavalid;                                           // mm_interconnect_0:cpu_0_instruction_master_readdatavalid -> cpu_0:i_readdatavalid
	wire  [31:0] cpu_3_data_master_readdata;                                                       // mm_interconnect_0:cpu_3_data_master_readdata -> cpu_3:d_readdata
	wire         cpu_3_data_master_waitrequest;                                                    // mm_interconnect_0:cpu_3_data_master_waitrequest -> cpu_3:d_waitrequest
	wire         cpu_3_data_master_debugaccess;                                                    // cpu_3:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_3_data_master_debugaccess
	wire  [21:0] cpu_3_data_master_address;                                                        // cpu_3:d_address -> mm_interconnect_0:cpu_3_data_master_address
	wire   [3:0] cpu_3_data_master_byteenable;                                                     // cpu_3:d_byteenable -> mm_interconnect_0:cpu_3_data_master_byteenable
	wire         cpu_3_data_master_read;                                                           // cpu_3:d_read -> mm_interconnect_0:cpu_3_data_master_read
	wire         cpu_3_data_master_readdatavalid;                                                  // mm_interconnect_0:cpu_3_data_master_readdatavalid -> cpu_3:d_readdatavalid
	wire         cpu_3_data_master_write;                                                          // cpu_3:d_write -> mm_interconnect_0:cpu_3_data_master_write
	wire  [31:0] cpu_3_data_master_writedata;                                                      // cpu_3:d_writedata -> mm_interconnect_0:cpu_3_data_master_writedata
	wire  [31:0] cpu_2_data_master_readdata;                                                       // mm_interconnect_0:cpu_2_data_master_readdata -> cpu_2:d_readdata
	wire         cpu_2_data_master_waitrequest;                                                    // mm_interconnect_0:cpu_2_data_master_waitrequest -> cpu_2:d_waitrequest
	wire         cpu_2_data_master_debugaccess;                                                    // cpu_2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_2_data_master_debugaccess
	wire  [21:0] cpu_2_data_master_address;                                                        // cpu_2:d_address -> mm_interconnect_0:cpu_2_data_master_address
	wire   [3:0] cpu_2_data_master_byteenable;                                                     // cpu_2:d_byteenable -> mm_interconnect_0:cpu_2_data_master_byteenable
	wire         cpu_2_data_master_read;                                                           // cpu_2:d_read -> mm_interconnect_0:cpu_2_data_master_read
	wire         cpu_2_data_master_readdatavalid;                                                  // mm_interconnect_0:cpu_2_data_master_readdatavalid -> cpu_2:d_readdatavalid
	wire         cpu_2_data_master_write;                                                          // cpu_2:d_write -> mm_interconnect_0:cpu_2_data_master_write
	wire  [31:0] cpu_2_data_master_writedata;                                                      // cpu_2:d_writedata -> mm_interconnect_0:cpu_2_data_master_writedata
	wire  [31:0] cpu_1_data_master_readdata;                                                       // mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	wire         cpu_1_data_master_waitrequest;                                                    // mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	wire         cpu_1_data_master_debugaccess;                                                    // cpu_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	wire  [21:0] cpu_1_data_master_address;                                                        // cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	wire   [3:0] cpu_1_data_master_byteenable;                                                     // cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	wire         cpu_1_data_master_read;                                                           // cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	wire         cpu_1_data_master_readdatavalid;                                                  // mm_interconnect_0:cpu_1_data_master_readdatavalid -> cpu_1:d_readdatavalid
	wire         cpu_1_data_master_write;                                                          // cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	wire  [31:0] cpu_1_data_master_writedata;                                                      // cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	wire  [31:0] cpu_3_instruction_master_readdata;                                                // mm_interconnect_0:cpu_3_instruction_master_readdata -> cpu_3:i_readdata
	wire         cpu_3_instruction_master_waitrequest;                                             // mm_interconnect_0:cpu_3_instruction_master_waitrequest -> cpu_3:i_waitrequest
	wire  [21:0] cpu_3_instruction_master_address;                                                 // cpu_3:i_address -> mm_interconnect_0:cpu_3_instruction_master_address
	wire         cpu_3_instruction_master_read;                                                    // cpu_3:i_read -> mm_interconnect_0:cpu_3_instruction_master_read
	wire         cpu_3_instruction_master_readdatavalid;                                           // mm_interconnect_0:cpu_3_instruction_master_readdatavalid -> cpu_3:i_readdatavalid
	wire  [31:0] cpu_2_instruction_master_readdata;                                                // mm_interconnect_0:cpu_2_instruction_master_readdata -> cpu_2:i_readdata
	wire         cpu_2_instruction_master_waitrequest;                                             // mm_interconnect_0:cpu_2_instruction_master_waitrequest -> cpu_2:i_waitrequest
	wire  [21:0] cpu_2_instruction_master_address;                                                 // cpu_2:i_address -> mm_interconnect_0:cpu_2_instruction_master_address
	wire         cpu_2_instruction_master_read;                                                    // cpu_2:i_read -> mm_interconnect_0:cpu_2_instruction_master_read
	wire         cpu_2_instruction_master_readdatavalid;                                           // mm_interconnect_0:cpu_2_instruction_master_readdatavalid -> cpu_2:i_readdatavalid
	wire  [31:0] cpu_1_instruction_master_readdata;                                                // mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	wire         cpu_1_instruction_master_waitrequest;                                             // mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	wire  [21:0] cpu_1_instruction_master_address;                                                 // cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	wire         cpu_1_instruction_master_read;                                                    // cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	wire         cpu_1_instruction_master_readdatavalid;                                           // mm_interconnect_0:cpu_1_instruction_master_readdatavalid -> cpu_1:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                           // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                        // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_hypervisor_debug_mem_slave_readdata;                            // hypervisor:debug_mem_slave_readdata -> mm_interconnect_0:hypervisor_debug_mem_slave_readdata
	wire         mm_interconnect_0_hypervisor_debug_mem_slave_waitrequest;                         // hypervisor:debug_mem_slave_waitrequest -> mm_interconnect_0:hypervisor_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_hypervisor_debug_mem_slave_debugaccess;                         // mm_interconnect_0:hypervisor_debug_mem_slave_debugaccess -> hypervisor:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_hypervisor_debug_mem_slave_address;                             // mm_interconnect_0:hypervisor_debug_mem_slave_address -> hypervisor:debug_mem_slave_address
	wire         mm_interconnect_0_hypervisor_debug_mem_slave_read;                                // mm_interconnect_0:hypervisor_debug_mem_slave_read -> hypervisor:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_hypervisor_debug_mem_slave_byteenable;                          // mm_interconnect_0:hypervisor_debug_mem_slave_byteenable -> hypervisor:debug_mem_slave_byteenable
	wire         mm_interconnect_0_hypervisor_debug_mem_slave_write;                               // mm_interconnect_0:hypervisor_debug_mem_slave_write -> hypervisor:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_hypervisor_debug_mem_slave_writedata;                           // mm_interconnect_0:hypervisor_debug_mem_slave_writedata -> hypervisor:debug_mem_slave_writedata
	wire         mm_interconnect_0_uart_rs_s1_chipselect;                                          // mm_interconnect_0:uart_rs_s1_chipselect -> uart_rs:chipselect
	wire  [15:0] mm_interconnect_0_uart_rs_s1_readdata;                                            // uart_rs:readdata -> mm_interconnect_0:uart_rs_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_rs_s1_address;                                             // mm_interconnect_0:uart_rs_s1_address -> uart_rs:address
	wire         mm_interconnect_0_uart_rs_s1_read;                                                // mm_interconnect_0:uart_rs_s1_read -> uart_rs:read_n
	wire         mm_interconnect_0_uart_rs_s1_begintransfer;                                       // mm_interconnect_0:uart_rs_s1_begintransfer -> uart_rs:begintransfer
	wire         mm_interconnect_0_uart_rs_s1_write;                                               // mm_interconnect_0:uart_rs_s1_write -> uart_rs:write_n
	wire  [15:0] mm_interconnect_0_uart_rs_s1_writedata;                                           // mm_interconnect_0:uart_rs_s1_writedata -> uart_rs:writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                                              // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                                                // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [15:0] mm_interconnect_0_ram_s1_address;                                                 // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                                              // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                                                   // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                                               // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                                                   // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire  [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_readdata;                                 // cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest;                              // cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess;                              // mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_0_debug_mem_slave_address;                                  // mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_read;                                     // mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_0_debug_mem_slave_byteenable;                               // mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_write;                                    // mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_writedata;                                // mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_cpu_1_debug_mem_slave_readdata;                                 // cpu_1:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest;                              // cpu_1:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess;                              // mm_interconnect_0:cpu_1_debug_mem_slave_debugaccess -> cpu_1:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_1_debug_mem_slave_address;                                  // mm_interconnect_0:cpu_1_debug_mem_slave_address -> cpu_1:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_read;                                     // mm_interconnect_0:cpu_1_debug_mem_slave_read -> cpu_1:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_1_debug_mem_slave_byteenable;                               // mm_interconnect_0:cpu_1_debug_mem_slave_byteenable -> cpu_1:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_1_debug_mem_slave_write;                                    // mm_interconnect_0:cpu_1_debug_mem_slave_write -> cpu_1:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_1_debug_mem_slave_writedata;                                // mm_interconnect_0:cpu_1_debug_mem_slave_writedata -> cpu_1:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_cpu_2_debug_mem_slave_readdata;                                 // cpu_2:debug_mem_slave_readdata -> mm_interconnect_0:cpu_2_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest;                              // cpu_2:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess;                              // mm_interconnect_0:cpu_2_debug_mem_slave_debugaccess -> cpu_2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_2_debug_mem_slave_address;                                  // mm_interconnect_0:cpu_2_debug_mem_slave_address -> cpu_2:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_2_debug_mem_slave_read;                                     // mm_interconnect_0:cpu_2_debug_mem_slave_read -> cpu_2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_2_debug_mem_slave_byteenable;                               // mm_interconnect_0:cpu_2_debug_mem_slave_byteenable -> cpu_2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_2_debug_mem_slave_write;                                    // mm_interconnect_0:cpu_2_debug_mem_slave_write -> cpu_2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_2_debug_mem_slave_writedata;                                // mm_interconnect_0:cpu_2_debug_mem_slave_writedata -> cpu_2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_cpu_3_debug_mem_slave_readdata;                                 // cpu_3:debug_mem_slave_readdata -> mm_interconnect_0:cpu_3_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_3_debug_mem_slave_waitrequest;                              // cpu_3:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_3_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_3_debug_mem_slave_debugaccess;                              // mm_interconnect_0:cpu_3_debug_mem_slave_debugaccess -> cpu_3:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_3_debug_mem_slave_address;                                  // mm_interconnect_0:cpu_3_debug_mem_slave_address -> cpu_3:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_3_debug_mem_slave_read;                                     // mm_interconnect_0:cpu_3_debug_mem_slave_read -> cpu_3:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_3_debug_mem_slave_byteenable;                               // mm_interconnect_0:cpu_3_debug_mem_slave_byteenable -> cpu_3:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_3_debug_mem_slave_write;                                    // mm_interconnect_0:cpu_3_debug_mem_slave_write -> cpu_3:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_3_debug_mem_slave_writedata;                                // mm_interconnect_0:cpu_3_debug_mem_slave_writedata -> cpu_3:debug_mem_slave_writedata
	wire  [31:0] cpu_0_irq_irq;                                                                    // irq_mapper:sender_irq -> cpu_0:irq
	wire  [31:0] cpu_1_irq_irq;                                                                    // irq_mapper_001:sender_irq -> cpu_1:irq
	wire  [31:0] cpu_2_irq_irq;                                                                    // irq_mapper_002:sender_irq -> cpu_2:irq
	wire  [31:0] cpu_3_irq_irq;                                                                    // irq_mapper_003:sender_irq -> cpu_3:irq
	wire         irq_mapper_004_receiver0_irq;                                                     // uart_rs:irq -> irq_mapper_004:receiver0_irq
	wire  [31:0] hypervisor_irq_irq;                                                               // irq_mapper_004:sender_irq -> hypervisor:irq
	wire         irq_mapper_receiver0_irq;                                                         // jtag_uart:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_004:receiver1_irq]
	wire         rst_controller_reset_out_reset;                                                   // rst_controller:reset_out -> [RAM:reset, cpu_0:reset_n, cpu_1:reset_n, cpu_2:reset_n, cpu_3:reset_n, hypervisor:reset_n, irq_mapper:reset, irq_mapper_001:reset, irq_mapper_002:reset, irq_mapper_003:reset, irq_mapper_004:reset, jtag_uart:rst_n, mm_interconnect_0:hypervisor_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, uart_rs:reset_n]
	wire         rst_controller_reset_out_reset_req;                                               // rst_controller:reset_req -> [RAM:reset_req, cpu_0:reset_req, cpu_1:reset_req, cpu_2:reset_req, cpu_3:reset_req, hypervisor:reset_req, rst_translator:reset_req_in]

	parallel_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	parallel_cpu_0 cpu_0 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (cpu_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_0_data_master_read),                              //                          .read
		.d_readdata                          (cpu_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_0_data_master_write),                             //                          .write
		.d_writedata                         (cpu_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_0_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                    //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (cpu_0_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (cpu_0_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (cpu_0_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (cpu_0_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (cpu_0_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (cpu_0_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (cpu_0_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (cpu_0_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (cpu_0_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (cpu_0_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (cpu_0_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (cpu_0_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (cpu_0_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (cpu_0_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (cpu_0_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (cpu_0_custom_instruction_master_multi_writerc),       //                          .multi_writerc
		.E_ci_combo_result                   (cpu_0_custom_instruction_master_result),              //                          .result
		.E_ci_combo_a                        (cpu_0_custom_instruction_master_a),                   //                          .a
		.E_ci_combo_b                        (cpu_0_custom_instruction_master_b),                   //                          .b
		.E_ci_combo_c                        (cpu_0_custom_instruction_master_c),                   //                          .c
		.E_ci_combo_dataa                    (cpu_0_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_combo_datab                    (cpu_0_custom_instruction_master_datab),               //                          .datab
		.E_ci_combo_estatus                  (cpu_0_custom_instruction_master_estatus),             //                          .estatus
		.E_ci_combo_ipending                 (cpu_0_custom_instruction_master_ipending),            //                          .ipending
		.E_ci_combo_n                        (cpu_0_custom_instruction_master_n),                   //                          .n
		.E_ci_combo_readra                   (cpu_0_custom_instruction_master_readra),              //                          .readra
		.E_ci_combo_readrb                   (cpu_0_custom_instruction_master_readrb),              //                          .readrb
		.E_ci_combo_writerc                  (cpu_0_custom_instruction_master_writerc)              //                          .writerc
	);

	parallel_cpu_1 cpu_1 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (cpu_1_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_1_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_1_data_master_read),                              //                          .read
		.d_readdata                          (cpu_1_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_1_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_1_data_master_write),                             //                          .write
		.d_writedata                         (cpu_1_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_1_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_1_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_1_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_1_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_1_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_1_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_1_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_1_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                    //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_1_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_1_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_1_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_1_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_1_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_1_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	parallel_cpu_2 cpu_2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (cpu_2_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_2_data_master_read),                              //                          .read
		.d_readdata                          (cpu_2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_2_data_master_write),                             //                          .write
		.d_writedata                         (cpu_2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_2_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                    //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_2_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (cpu_2_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (cpu_2_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (cpu_2_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (cpu_2_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (cpu_2_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (cpu_2_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (cpu_2_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (cpu_2_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (cpu_2_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (cpu_2_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (cpu_2_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (cpu_2_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (cpu_2_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (cpu_2_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (cpu_2_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (cpu_2_custom_instruction_master_multi_writerc),       //                          .multi_writerc
		.E_ci_combo_result                   (cpu_2_custom_instruction_master_result),              //                          .result
		.E_ci_combo_a                        (cpu_2_custom_instruction_master_a),                   //                          .a
		.E_ci_combo_b                        (cpu_2_custom_instruction_master_b),                   //                          .b
		.E_ci_combo_c                        (cpu_2_custom_instruction_master_c),                   //                          .c
		.E_ci_combo_dataa                    (cpu_2_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_combo_datab                    (cpu_2_custom_instruction_master_datab),               //                          .datab
		.E_ci_combo_estatus                  (cpu_2_custom_instruction_master_estatus),             //                          .estatus
		.E_ci_combo_ipending                 (cpu_2_custom_instruction_master_ipending),            //                          .ipending
		.E_ci_combo_n                        (cpu_2_custom_instruction_master_n),                   //                          .n
		.E_ci_combo_readra                   (cpu_2_custom_instruction_master_readra),              //                          .readra
		.E_ci_combo_readrb                   (cpu_2_custom_instruction_master_readrb),              //                          .readrb
		.E_ci_combo_writerc                  (cpu_2_custom_instruction_master_writerc)              //                          .writerc
	);

	parallel_cpu_3 cpu_3 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (cpu_3_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_3_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_3_data_master_read),                              //                          .read
		.d_readdata                          (cpu_3_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_3_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_3_data_master_write),                             //                          .write
		.d_writedata                         (cpu_3_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_3_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_3_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_3_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_3_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_3_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_3_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_3_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_3_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                    //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_3_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_3_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_3_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_3_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_3_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_3_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_3_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_3_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (cpu_3_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (cpu_3_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (cpu_3_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (cpu_3_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (cpu_3_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (cpu_3_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (cpu_3_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (cpu_3_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (cpu_3_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (cpu_3_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (cpu_3_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (cpu_3_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (cpu_3_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (cpu_3_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (cpu_3_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (cpu_3_custom_instruction_master_multi_writerc),       //                          .multi_writerc
		.E_ci_combo_result                   (cpu_3_custom_instruction_master_result),              //                          .result
		.E_ci_combo_a                        (cpu_3_custom_instruction_master_a),                   //                          .a
		.E_ci_combo_b                        (cpu_3_custom_instruction_master_b),                   //                          .b
		.E_ci_combo_c                        (cpu_3_custom_instruction_master_c),                   //                          .c
		.E_ci_combo_dataa                    (cpu_3_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_combo_datab                    (cpu_3_custom_instruction_master_datab),               //                          .datab
		.E_ci_combo_estatus                  (cpu_3_custom_instruction_master_estatus),             //                          .estatus
		.E_ci_combo_ipending                 (cpu_3_custom_instruction_master_ipending),            //                          .ipending
		.E_ci_combo_n                        (cpu_3_custom_instruction_master_n),                   //                          .n
		.E_ci_combo_readra                   (cpu_3_custom_instruction_master_readra),              //                          .readra
		.E_ci_combo_readrb                   (cpu_3_custom_instruction_master_readrb),              //                          .readrb
		.E_ci_combo_writerc                  (cpu_3_custom_instruction_master_writerc)              //                          .writerc
	);

	parallel_fpu_0 #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1),
		.comparison_present (1)
	) fpu_0 (
		.s1_dataa     (cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	parallel_fpu_0 #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1),
		.comparison_present (1)
	) fpu_1 (
		.s1_dataa     (), // s1.dataa
		.s1_datab     (), //   .datab
		.s1_n         (), //   .n
		.s1_result    (), //   .result
		.s2_clk       (), // s2.clk
		.s2_clk_en    (), //   .clk_en
		.s2_dataa     (), //   .dataa
		.s2_datab     (), //   .datab
		.s2_n         (), //   .n
		.s2_reset     (), //   .reset
		.s2_reset_req (), //   .reset_req
		.s2_start     (), //   .start
		.s2_done      (), //   .done
		.s2_result    ()  //   .result
	);

	parallel_fpu_0 #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1),
		.comparison_present (1)
	) fpu_2 (
		.s1_dataa     (cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	parallel_fpu_0 #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1),
		.comparison_present (1)
	) fpu_3 (
		.s1_dataa     (cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	parallel_hypervisor hypervisor (
		.clk                                 (clk_clk),                                                  //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                          //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                       //                          .reset_req
		.d_address                           (hypervisor_data_master_address),                           //               data_master.address
		.d_byteenable                        (hypervisor_data_master_byteenable),                        //                          .byteenable
		.d_read                              (hypervisor_data_master_read),                              //                          .read
		.d_readdata                          (hypervisor_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (hypervisor_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (hypervisor_data_master_write),                             //                          .write
		.d_writedata                         (hypervisor_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (hypervisor_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (hypervisor_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (hypervisor_instruction_master_address),                    //        instruction_master.address
		.i_read                              (hypervisor_instruction_master_read),                       //                          .read
		.i_readdata                          (hypervisor_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (hypervisor_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (hypervisor_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (hypervisor_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (hypervisor_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_hypervisor_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_hypervisor_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_hypervisor_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_hypervisor_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_hypervisor_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_hypervisor_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_hypervisor_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_hypervisor_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (hypervisor_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (hypervisor_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (hypervisor_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (hypervisor_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (hypervisor_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (hypervisor_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (hypervisor_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (hypervisor_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (hypervisor_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (hypervisor_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (hypervisor_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (hypervisor_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (hypervisor_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (hypervisor_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (hypervisor_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (hypervisor_custom_instruction_master_multi_writerc),       //                          .multi_writerc
		.E_ci_combo_result                   (hypervisor_custom_instruction_master_result),              //                          .result
		.E_ci_combo_a                        (hypervisor_custom_instruction_master_a),                   //                          .a
		.E_ci_combo_b                        (hypervisor_custom_instruction_master_b),                   //                          .b
		.E_ci_combo_c                        (hypervisor_custom_instruction_master_c),                   //                          .c
		.E_ci_combo_dataa                    (hypervisor_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_combo_datab                    (hypervisor_custom_instruction_master_datab),               //                          .datab
		.E_ci_combo_estatus                  (hypervisor_custom_instruction_master_estatus),             //                          .estatus
		.E_ci_combo_ipending                 (hypervisor_custom_instruction_master_ipending),            //                          .ipending
		.E_ci_combo_n                        (hypervisor_custom_instruction_master_n),                   //                          .n
		.E_ci_combo_readra                   (hypervisor_custom_instruction_master_readra),              //                          .readra
		.E_ci_combo_readrb                   (hypervisor_custom_instruction_master_readrb),              //                          .readrb
		.E_ci_combo_writerc                  (hypervisor_custom_instruction_master_writerc)              //                          .writerc
	);

	parallel_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	parallel_fpu_0 #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1),
		.comparison_present (1)
	) nios2_fpu (
		.s1_dataa     (hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	parallel_uart_rs uart_rs (
		.clk           (clk_clk),                                    //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address       (mm_interconnect_0_uart_rs_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_rs_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_rs_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_rs_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_rs_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_rs_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_rs_s1_readdata),      //                    .readdata
		.rxd           (uart_0_external_connection_rxd),             // external_connection.export
		.txd           (uart_0_external_connection_txd),             //                    .export
		.irq           (irq_mapper_004_receiver0_irq)                //                 irq.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) hypervisor_custom_instruction_master_translator (
		.ci_slave_dataa            (hypervisor_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (hypervisor_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (hypervisor_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (hypervisor_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (hypervisor_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (hypervisor_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (hypervisor_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (hypervisor_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (hypervisor_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (hypervisor_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (hypervisor_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (hypervisor_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (hypervisor_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (hypervisor_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (hypervisor_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (hypervisor_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (hypervisor_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (hypervisor_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (hypervisor_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (hypervisor_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (hypervisor_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (hypervisor_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (hypervisor_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (hypervisor_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (hypervisor_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (hypervisor_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (hypervisor_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (hypervisor_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (hypervisor_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (hypervisor_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (hypervisor_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (hypervisor_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (hypervisor_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (hypervisor_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (hypervisor_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (hypervisor_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (hypervisor_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (hypervisor_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (hypervisor_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (hypervisor_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (hypervisor_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (hypervisor_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (hypervisor_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (hypervisor_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (hypervisor_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (hypervisor_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (hypervisor_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (hypervisor_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (hypervisor_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (hypervisor_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (hypervisor_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (hypervisor_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (hypervisor_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (hypervisor_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (hypervisor_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (hypervisor_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	parallel_hypervisor_custom_instruction_master_comb_xconnect hypervisor_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (hypervisor_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (hypervisor_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (hypervisor_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (hypervisor_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (hypervisor_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (hypervisor_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (hypervisor_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (hypervisor_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (hypervisor_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (hypervisor_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (hypervisor_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (hypervisor_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) hypervisor_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (hypervisor_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (hypervisor_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                             // (terminated)
		.ci_master_readrb    (),                                                                             // (terminated)
		.ci_master_writerc   (),                                                                             // (terminated)
		.ci_master_a         (),                                                                             // (terminated)
		.ci_master_b         (),                                                                             // (terminated)
		.ci_master_c         (),                                                                             // (terminated)
		.ci_master_ipending  (),                                                                             // (terminated)
		.ci_master_estatus   (),                                                                             // (terminated)
		.ci_master_clk       (),                                                                             // (terminated)
		.ci_master_clken     (),                                                                             // (terminated)
		.ci_master_reset_req (),                                                                             // (terminated)
		.ci_master_reset     (),                                                                             // (terminated)
		.ci_master_start     (),                                                                             // (terminated)
		.ci_master_done      (1'b0),                                                                         // (terminated)
		.ci_slave_clk        (1'b0),                                                                         // (terminated)
		.ci_slave_clken      (1'b0),                                                                         // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                         // (terminated)
		.ci_slave_reset      (1'b0),                                                                         // (terminated)
		.ci_slave_start      (1'b0),                                                                         // (terminated)
		.ci_slave_done       ()                                                                              // (terminated)
	);

	parallel_hypervisor_custom_instruction_master_multi_xconnect hypervisor_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (hypervisor_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (hypervisor_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (hypervisor_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (hypervisor_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (hypervisor_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (hypervisor_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (hypervisor_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (hypervisor_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (hypervisor_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (hypervisor_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                          //           .ipending
		.ci_slave_estatus     (),                                                                          //           .estatus
		.ci_slave_clk         (hypervisor_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (hypervisor_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (hypervisor_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (hypervisor_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (hypervisor_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (hypervisor_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) hypervisor_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (hypervisor_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (hypervisor_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                                 // (terminated)
		.ci_master_readrb    (),                                                                                 // (terminated)
		.ci_master_writerc   (),                                                                                 // (terminated)
		.ci_master_a         (),                                                                                 // (terminated)
		.ci_master_b         (),                                                                                 // (terminated)
		.ci_master_c         (),                                                                                 // (terminated)
		.ci_master_ipending  (),                                                                                 // (terminated)
		.ci_master_estatus   ()                                                                                  // (terminated)
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) cpu_2_custom_instruction_master_translator (
		.ci_slave_dataa            (cpu_2_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (cpu_2_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (cpu_2_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (cpu_2_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (cpu_2_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (cpu_2_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (cpu_2_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (cpu_2_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (cpu_2_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (cpu_2_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (cpu_2_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (cpu_2_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (cpu_2_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (cpu_2_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (cpu_2_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (cpu_2_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (cpu_2_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (cpu_2_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (cpu_2_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (cpu_2_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (cpu_2_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (cpu_2_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (cpu_2_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (cpu_2_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (cpu_2_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (cpu_2_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (cpu_2_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (cpu_2_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (cpu_2_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (cpu_2_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (cpu_2_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (cpu_2_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (cpu_2_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (cpu_2_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (cpu_2_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (cpu_2_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (cpu_2_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (cpu_2_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (cpu_2_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (cpu_2_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (cpu_2_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (cpu_2_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (cpu_2_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (cpu_2_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (cpu_2_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (cpu_2_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (cpu_2_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (cpu_2_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (cpu_2_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (cpu_2_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (cpu_2_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (cpu_2_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (cpu_2_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (cpu_2_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (cpu_2_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (cpu_2_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	parallel_hypervisor_custom_instruction_master_comb_xconnect cpu_2_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (cpu_2_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (cpu_2_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (cpu_2_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (cpu_2_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (cpu_2_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (cpu_2_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (cpu_2_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (cpu_2_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (cpu_2_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (cpu_2_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (cpu_2_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (cpu_2_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) cpu_2_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (cpu_2_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (cpu_2_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_clk       (),                                                                        // (terminated)
		.ci_master_clken     (),                                                                        // (terminated)
		.ci_master_reset_req (),                                                                        // (terminated)
		.ci_master_reset     (),                                                                        // (terminated)
		.ci_master_start     (),                                                                        // (terminated)
		.ci_master_done      (1'b0),                                                                    // (terminated)
		.ci_slave_clk        (1'b0),                                                                    // (terminated)
		.ci_slave_clken      (1'b0),                                                                    // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                    // (terminated)
		.ci_slave_reset      (1'b0),                                                                    // (terminated)
		.ci_slave_start      (1'b0),                                                                    // (terminated)
		.ci_slave_done       ()                                                                         // (terminated)
	);

	parallel_hypervisor_custom_instruction_master_multi_xconnect cpu_2_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (cpu_2_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (cpu_2_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (cpu_2_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (cpu_2_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (cpu_2_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (cpu_2_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (cpu_2_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (cpu_2_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (cpu_2_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (cpu_2_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                     //           .ipending
		.ci_slave_estatus     (),                                                                     //           .estatus
		.ci_slave_clk         (cpu_2_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (cpu_2_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (cpu_2_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (cpu_2_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (cpu_2_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (cpu_2_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) cpu_2_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (cpu_2_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (cpu_2_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                            // (terminated)
		.ci_master_readrb    (),                                                                            // (terminated)
		.ci_master_writerc   (),                                                                            // (terminated)
		.ci_master_a         (),                                                                            // (terminated)
		.ci_master_b         (),                                                                            // (terminated)
		.ci_master_c         (),                                                                            // (terminated)
		.ci_master_ipending  (),                                                                            // (terminated)
		.ci_master_estatus   ()                                                                             // (terminated)
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) cpu_3_custom_instruction_master_translator (
		.ci_slave_dataa            (cpu_3_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (cpu_3_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (cpu_3_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (cpu_3_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (cpu_3_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (cpu_3_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (cpu_3_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (cpu_3_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (cpu_3_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (cpu_3_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (cpu_3_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (cpu_3_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (cpu_3_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (cpu_3_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (cpu_3_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (cpu_3_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (cpu_3_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (cpu_3_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (cpu_3_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (cpu_3_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (cpu_3_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (cpu_3_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (cpu_3_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (cpu_3_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (cpu_3_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (cpu_3_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (cpu_3_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (cpu_3_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (cpu_3_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (cpu_3_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (cpu_3_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (cpu_3_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (cpu_3_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (cpu_3_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (cpu_3_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (cpu_3_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (cpu_3_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (cpu_3_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (cpu_3_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (cpu_3_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (cpu_3_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (cpu_3_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (cpu_3_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (cpu_3_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (cpu_3_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (cpu_3_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (cpu_3_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (cpu_3_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (cpu_3_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (cpu_3_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (cpu_3_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (cpu_3_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (cpu_3_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (cpu_3_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (cpu_3_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (cpu_3_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	parallel_hypervisor_custom_instruction_master_comb_xconnect cpu_3_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (cpu_3_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (cpu_3_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (cpu_3_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (cpu_3_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (cpu_3_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (cpu_3_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (cpu_3_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (cpu_3_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (cpu_3_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (cpu_3_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (cpu_3_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (cpu_3_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) cpu_3_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (cpu_3_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (cpu_3_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_clk       (),                                                                        // (terminated)
		.ci_master_clken     (),                                                                        // (terminated)
		.ci_master_reset_req (),                                                                        // (terminated)
		.ci_master_reset     (),                                                                        // (terminated)
		.ci_master_start     (),                                                                        // (terminated)
		.ci_master_done      (1'b0),                                                                    // (terminated)
		.ci_slave_clk        (1'b0),                                                                    // (terminated)
		.ci_slave_clken      (1'b0),                                                                    // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                    // (terminated)
		.ci_slave_reset      (1'b0),                                                                    // (terminated)
		.ci_slave_start      (1'b0),                                                                    // (terminated)
		.ci_slave_done       ()                                                                         // (terminated)
	);

	parallel_hypervisor_custom_instruction_master_multi_xconnect cpu_3_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (cpu_3_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (cpu_3_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (cpu_3_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (cpu_3_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (cpu_3_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (cpu_3_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (cpu_3_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (cpu_3_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (cpu_3_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (cpu_3_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                     //           .ipending
		.ci_slave_estatus     (),                                                                     //           .estatus
		.ci_slave_clk         (cpu_3_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (cpu_3_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (cpu_3_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (cpu_3_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (cpu_3_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (cpu_3_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) cpu_3_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (cpu_3_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (cpu_3_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                            // (terminated)
		.ci_master_readrb    (),                                                                            // (terminated)
		.ci_master_writerc   (),                                                                            // (terminated)
		.ci_master_a         (),                                                                            // (terminated)
		.ci_master_b         (),                                                                            // (terminated)
		.ci_master_c         (),                                                                            // (terminated)
		.ci_master_ipending  (),                                                                            // (terminated)
		.ci_master_estatus   ()                                                                             // (terminated)
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) cpu_0_custom_instruction_master_translator (
		.ci_slave_dataa            (cpu_0_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (cpu_0_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (cpu_0_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (cpu_0_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (cpu_0_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (cpu_0_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (cpu_0_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (cpu_0_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (cpu_0_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (cpu_0_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (cpu_0_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (cpu_0_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (cpu_0_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (cpu_0_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (cpu_0_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (cpu_0_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (cpu_0_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (cpu_0_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (cpu_0_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (cpu_0_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (cpu_0_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (cpu_0_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (cpu_0_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (cpu_0_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (cpu_0_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (cpu_0_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (cpu_0_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (cpu_0_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (cpu_0_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (cpu_0_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (cpu_0_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (cpu_0_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (cpu_0_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (cpu_0_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (cpu_0_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (cpu_0_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (cpu_0_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (cpu_0_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (cpu_0_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (cpu_0_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (cpu_0_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (cpu_0_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (cpu_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (cpu_0_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (cpu_0_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (cpu_0_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (cpu_0_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (cpu_0_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (cpu_0_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (cpu_0_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (cpu_0_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (cpu_0_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (cpu_0_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (cpu_0_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (cpu_0_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (cpu_0_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	parallel_hypervisor_custom_instruction_master_comb_xconnect cpu_0_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (cpu_0_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (cpu_0_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (cpu_0_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (cpu_0_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (cpu_0_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (cpu_0_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (cpu_0_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (cpu_0_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (cpu_0_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (cpu_0_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (cpu_0_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (cpu_0_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) cpu_0_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (cpu_0_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (cpu_0_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_clk       (),                                                                        // (terminated)
		.ci_master_clken     (),                                                                        // (terminated)
		.ci_master_reset_req (),                                                                        // (terminated)
		.ci_master_reset     (),                                                                        // (terminated)
		.ci_master_start     (),                                                                        // (terminated)
		.ci_master_done      (1'b0),                                                                    // (terminated)
		.ci_slave_clk        (1'b0),                                                                    // (terminated)
		.ci_slave_clken      (1'b0),                                                                    // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                    // (terminated)
		.ci_slave_reset      (1'b0),                                                                    // (terminated)
		.ci_slave_start      (1'b0),                                                                    // (terminated)
		.ci_slave_done       ()                                                                         // (terminated)
	);

	parallel_hypervisor_custom_instruction_master_multi_xconnect cpu_0_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (cpu_0_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (cpu_0_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (cpu_0_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (cpu_0_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (cpu_0_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (cpu_0_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (cpu_0_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (cpu_0_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (cpu_0_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (cpu_0_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                     //           .ipending
		.ci_slave_estatus     (),                                                                     //           .estatus
		.ci_slave_clk         (cpu_0_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (cpu_0_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (cpu_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (cpu_0_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (cpu_0_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (cpu_0_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) cpu_0_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (cpu_0_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (cpu_0_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                            // (terminated)
		.ci_master_readrb    (),                                                                            // (terminated)
		.ci_master_writerc   (),                                                                            // (terminated)
		.ci_master_a         (),                                                                            // (terminated)
		.ci_master_b         (),                                                                            // (terminated)
		.ci_master_c         (),                                                                            // (terminated)
		.ci_master_ipending  (),                                                                            // (terminated)
		.ci_master_estatus   ()                                                                             // (terminated)
	);

	parallel_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                (clk_clk),                                                   //                              clk_0_clk.clk
		.hypervisor_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // hypervisor_reset_reset_bridge_in_reset.reset
		.cpu_0_data_master_address                    (cpu_0_data_master_address),                                 //                      cpu_0_data_master.address
		.cpu_0_data_master_waitrequest                (cpu_0_data_master_waitrequest),                             //                                       .waitrequest
		.cpu_0_data_master_byteenable                 (cpu_0_data_master_byteenable),                              //                                       .byteenable
		.cpu_0_data_master_read                       (cpu_0_data_master_read),                                    //                                       .read
		.cpu_0_data_master_readdata                   (cpu_0_data_master_readdata),                                //                                       .readdata
		.cpu_0_data_master_readdatavalid              (cpu_0_data_master_readdatavalid),                           //                                       .readdatavalid
		.cpu_0_data_master_write                      (cpu_0_data_master_write),                                   //                                       .write
		.cpu_0_data_master_writedata                  (cpu_0_data_master_writedata),                               //                                       .writedata
		.cpu_0_data_master_debugaccess                (cpu_0_data_master_debugaccess),                             //                                       .debugaccess
		.cpu_0_instruction_master_address             (cpu_0_instruction_master_address),                          //               cpu_0_instruction_master.address
		.cpu_0_instruction_master_waitrequest         (cpu_0_instruction_master_waitrequest),                      //                                       .waitrequest
		.cpu_0_instruction_master_read                (cpu_0_instruction_master_read),                             //                                       .read
		.cpu_0_instruction_master_readdata            (cpu_0_instruction_master_readdata),                         //                                       .readdata
		.cpu_0_instruction_master_readdatavalid       (cpu_0_instruction_master_readdatavalid),                    //                                       .readdatavalid
		.cpu_1_data_master_address                    (cpu_1_data_master_address),                                 //                      cpu_1_data_master.address
		.cpu_1_data_master_waitrequest                (cpu_1_data_master_waitrequest),                             //                                       .waitrequest
		.cpu_1_data_master_byteenable                 (cpu_1_data_master_byteenable),                              //                                       .byteenable
		.cpu_1_data_master_read                       (cpu_1_data_master_read),                                    //                                       .read
		.cpu_1_data_master_readdata                   (cpu_1_data_master_readdata),                                //                                       .readdata
		.cpu_1_data_master_readdatavalid              (cpu_1_data_master_readdatavalid),                           //                                       .readdatavalid
		.cpu_1_data_master_write                      (cpu_1_data_master_write),                                   //                                       .write
		.cpu_1_data_master_writedata                  (cpu_1_data_master_writedata),                               //                                       .writedata
		.cpu_1_data_master_debugaccess                (cpu_1_data_master_debugaccess),                             //                                       .debugaccess
		.cpu_1_instruction_master_address             (cpu_1_instruction_master_address),                          //               cpu_1_instruction_master.address
		.cpu_1_instruction_master_waitrequest         (cpu_1_instruction_master_waitrequest),                      //                                       .waitrequest
		.cpu_1_instruction_master_read                (cpu_1_instruction_master_read),                             //                                       .read
		.cpu_1_instruction_master_readdata            (cpu_1_instruction_master_readdata),                         //                                       .readdata
		.cpu_1_instruction_master_readdatavalid       (cpu_1_instruction_master_readdatavalid),                    //                                       .readdatavalid
		.cpu_2_data_master_address                    (cpu_2_data_master_address),                                 //                      cpu_2_data_master.address
		.cpu_2_data_master_waitrequest                (cpu_2_data_master_waitrequest),                             //                                       .waitrequest
		.cpu_2_data_master_byteenable                 (cpu_2_data_master_byteenable),                              //                                       .byteenable
		.cpu_2_data_master_read                       (cpu_2_data_master_read),                                    //                                       .read
		.cpu_2_data_master_readdata                   (cpu_2_data_master_readdata),                                //                                       .readdata
		.cpu_2_data_master_readdatavalid              (cpu_2_data_master_readdatavalid),                           //                                       .readdatavalid
		.cpu_2_data_master_write                      (cpu_2_data_master_write),                                   //                                       .write
		.cpu_2_data_master_writedata                  (cpu_2_data_master_writedata),                               //                                       .writedata
		.cpu_2_data_master_debugaccess                (cpu_2_data_master_debugaccess),                             //                                       .debugaccess
		.cpu_2_instruction_master_address             (cpu_2_instruction_master_address),                          //               cpu_2_instruction_master.address
		.cpu_2_instruction_master_waitrequest         (cpu_2_instruction_master_waitrequest),                      //                                       .waitrequest
		.cpu_2_instruction_master_read                (cpu_2_instruction_master_read),                             //                                       .read
		.cpu_2_instruction_master_readdata            (cpu_2_instruction_master_readdata),                         //                                       .readdata
		.cpu_2_instruction_master_readdatavalid       (cpu_2_instruction_master_readdatavalid),                    //                                       .readdatavalid
		.cpu_3_data_master_address                    (cpu_3_data_master_address),                                 //                      cpu_3_data_master.address
		.cpu_3_data_master_waitrequest                (cpu_3_data_master_waitrequest),                             //                                       .waitrequest
		.cpu_3_data_master_byteenable                 (cpu_3_data_master_byteenable),                              //                                       .byteenable
		.cpu_3_data_master_read                       (cpu_3_data_master_read),                                    //                                       .read
		.cpu_3_data_master_readdata                   (cpu_3_data_master_readdata),                                //                                       .readdata
		.cpu_3_data_master_readdatavalid              (cpu_3_data_master_readdatavalid),                           //                                       .readdatavalid
		.cpu_3_data_master_write                      (cpu_3_data_master_write),                                   //                                       .write
		.cpu_3_data_master_writedata                  (cpu_3_data_master_writedata),                               //                                       .writedata
		.cpu_3_data_master_debugaccess                (cpu_3_data_master_debugaccess),                             //                                       .debugaccess
		.cpu_3_instruction_master_address             (cpu_3_instruction_master_address),                          //               cpu_3_instruction_master.address
		.cpu_3_instruction_master_waitrequest         (cpu_3_instruction_master_waitrequest),                      //                                       .waitrequest
		.cpu_3_instruction_master_read                (cpu_3_instruction_master_read),                             //                                       .read
		.cpu_3_instruction_master_readdata            (cpu_3_instruction_master_readdata),                         //                                       .readdata
		.cpu_3_instruction_master_readdatavalid       (cpu_3_instruction_master_readdatavalid),                    //                                       .readdatavalid
		.hypervisor_data_master_address               (hypervisor_data_master_address),                            //                 hypervisor_data_master.address
		.hypervisor_data_master_waitrequest           (hypervisor_data_master_waitrequest),                        //                                       .waitrequest
		.hypervisor_data_master_byteenable            (hypervisor_data_master_byteenable),                         //                                       .byteenable
		.hypervisor_data_master_read                  (hypervisor_data_master_read),                               //                                       .read
		.hypervisor_data_master_readdata              (hypervisor_data_master_readdata),                           //                                       .readdata
		.hypervisor_data_master_readdatavalid         (hypervisor_data_master_readdatavalid),                      //                                       .readdatavalid
		.hypervisor_data_master_write                 (hypervisor_data_master_write),                              //                                       .write
		.hypervisor_data_master_writedata             (hypervisor_data_master_writedata),                          //                                       .writedata
		.hypervisor_data_master_debugaccess           (hypervisor_data_master_debugaccess),                        //                                       .debugaccess
		.hypervisor_instruction_master_address        (hypervisor_instruction_master_address),                     //          hypervisor_instruction_master.address
		.hypervisor_instruction_master_waitrequest    (hypervisor_instruction_master_waitrequest),                 //                                       .waitrequest
		.hypervisor_instruction_master_read           (hypervisor_instruction_master_read),                        //                                       .read
		.hypervisor_instruction_master_readdata       (hypervisor_instruction_master_readdata),                    //                                       .readdata
		.hypervisor_instruction_master_readdatavalid  (hypervisor_instruction_master_readdatavalid),               //                                       .readdatavalid
		.cpu_0_debug_mem_slave_address                (mm_interconnect_0_cpu_0_debug_mem_slave_address),           //                  cpu_0_debug_mem_slave.address
		.cpu_0_debug_mem_slave_write                  (mm_interconnect_0_cpu_0_debug_mem_slave_write),             //                                       .write
		.cpu_0_debug_mem_slave_read                   (mm_interconnect_0_cpu_0_debug_mem_slave_read),              //                                       .read
		.cpu_0_debug_mem_slave_readdata               (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),          //                                       .readdata
		.cpu_0_debug_mem_slave_writedata              (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),         //                                       .writedata
		.cpu_0_debug_mem_slave_byteenable             (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),        //                                       .byteenable
		.cpu_0_debug_mem_slave_waitrequest            (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest),       //                                       .waitrequest
		.cpu_0_debug_mem_slave_debugaccess            (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess),       //                                       .debugaccess
		.cpu_1_debug_mem_slave_address                (mm_interconnect_0_cpu_1_debug_mem_slave_address),           //                  cpu_1_debug_mem_slave.address
		.cpu_1_debug_mem_slave_write                  (mm_interconnect_0_cpu_1_debug_mem_slave_write),             //                                       .write
		.cpu_1_debug_mem_slave_read                   (mm_interconnect_0_cpu_1_debug_mem_slave_read),              //                                       .read
		.cpu_1_debug_mem_slave_readdata               (mm_interconnect_0_cpu_1_debug_mem_slave_readdata),          //                                       .readdata
		.cpu_1_debug_mem_slave_writedata              (mm_interconnect_0_cpu_1_debug_mem_slave_writedata),         //                                       .writedata
		.cpu_1_debug_mem_slave_byteenable             (mm_interconnect_0_cpu_1_debug_mem_slave_byteenable),        //                                       .byteenable
		.cpu_1_debug_mem_slave_waitrequest            (mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest),       //                                       .waitrequest
		.cpu_1_debug_mem_slave_debugaccess            (mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess),       //                                       .debugaccess
		.cpu_2_debug_mem_slave_address                (mm_interconnect_0_cpu_2_debug_mem_slave_address),           //                  cpu_2_debug_mem_slave.address
		.cpu_2_debug_mem_slave_write                  (mm_interconnect_0_cpu_2_debug_mem_slave_write),             //                                       .write
		.cpu_2_debug_mem_slave_read                   (mm_interconnect_0_cpu_2_debug_mem_slave_read),              //                                       .read
		.cpu_2_debug_mem_slave_readdata               (mm_interconnect_0_cpu_2_debug_mem_slave_readdata),          //                                       .readdata
		.cpu_2_debug_mem_slave_writedata              (mm_interconnect_0_cpu_2_debug_mem_slave_writedata),         //                                       .writedata
		.cpu_2_debug_mem_slave_byteenable             (mm_interconnect_0_cpu_2_debug_mem_slave_byteenable),        //                                       .byteenable
		.cpu_2_debug_mem_slave_waitrequest            (mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest),       //                                       .waitrequest
		.cpu_2_debug_mem_slave_debugaccess            (mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess),       //                                       .debugaccess
		.cpu_3_debug_mem_slave_address                (mm_interconnect_0_cpu_3_debug_mem_slave_address),           //                  cpu_3_debug_mem_slave.address
		.cpu_3_debug_mem_slave_write                  (mm_interconnect_0_cpu_3_debug_mem_slave_write),             //                                       .write
		.cpu_3_debug_mem_slave_read                   (mm_interconnect_0_cpu_3_debug_mem_slave_read),              //                                       .read
		.cpu_3_debug_mem_slave_readdata               (mm_interconnect_0_cpu_3_debug_mem_slave_readdata),          //                                       .readdata
		.cpu_3_debug_mem_slave_writedata              (mm_interconnect_0_cpu_3_debug_mem_slave_writedata),         //                                       .writedata
		.cpu_3_debug_mem_slave_byteenable             (mm_interconnect_0_cpu_3_debug_mem_slave_byteenable),        //                                       .byteenable
		.cpu_3_debug_mem_slave_waitrequest            (mm_interconnect_0_cpu_3_debug_mem_slave_waitrequest),       //                                       .waitrequest
		.cpu_3_debug_mem_slave_debugaccess            (mm_interconnect_0_cpu_3_debug_mem_slave_debugaccess),       //                                       .debugaccess
		.hypervisor_debug_mem_slave_address           (mm_interconnect_0_hypervisor_debug_mem_slave_address),      //             hypervisor_debug_mem_slave.address
		.hypervisor_debug_mem_slave_write             (mm_interconnect_0_hypervisor_debug_mem_slave_write),        //                                       .write
		.hypervisor_debug_mem_slave_read              (mm_interconnect_0_hypervisor_debug_mem_slave_read),         //                                       .read
		.hypervisor_debug_mem_slave_readdata          (mm_interconnect_0_hypervisor_debug_mem_slave_readdata),     //                                       .readdata
		.hypervisor_debug_mem_slave_writedata         (mm_interconnect_0_hypervisor_debug_mem_slave_writedata),    //                                       .writedata
		.hypervisor_debug_mem_slave_byteenable        (mm_interconnect_0_hypervisor_debug_mem_slave_byteenable),   //                                       .byteenable
		.hypervisor_debug_mem_slave_waitrequest       (mm_interconnect_0_hypervisor_debug_mem_slave_waitrequest),  //                                       .waitrequest
		.hypervisor_debug_mem_slave_debugaccess       (mm_interconnect_0_hypervisor_debug_mem_slave_debugaccess),  //                                       .debugaccess
		.jtag_uart_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                       .write
		.jtag_uart_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                       .read
		.jtag_uart_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.RAM_s1_address                               (mm_interconnect_0_ram_s1_address),                          //                                 RAM_s1.address
		.RAM_s1_write                                 (mm_interconnect_0_ram_s1_write),                            //                                       .write
		.RAM_s1_readdata                              (mm_interconnect_0_ram_s1_readdata),                         //                                       .readdata
		.RAM_s1_writedata                             (mm_interconnect_0_ram_s1_writedata),                        //                                       .writedata
		.RAM_s1_byteenable                            (mm_interconnect_0_ram_s1_byteenable),                       //                                       .byteenable
		.RAM_s1_chipselect                            (mm_interconnect_0_ram_s1_chipselect),                       //                                       .chipselect
		.RAM_s1_clken                                 (mm_interconnect_0_ram_s1_clken),                            //                                       .clken
		.uart_rs_s1_address                           (mm_interconnect_0_uart_rs_s1_address),                      //                             uart_rs_s1.address
		.uart_rs_s1_write                             (mm_interconnect_0_uart_rs_s1_write),                        //                                       .write
		.uart_rs_s1_read                              (mm_interconnect_0_uart_rs_s1_read),                         //                                       .read
		.uart_rs_s1_readdata                          (mm_interconnect_0_uart_rs_s1_readdata),                     //                                       .readdata
		.uart_rs_s1_writedata                         (mm_interconnect_0_uart_rs_s1_writedata),                    //                                       .writedata
		.uart_rs_s1_begintransfer                     (mm_interconnect_0_uart_rs_s1_begintransfer),                //                                       .begintransfer
		.uart_rs_s1_chipselect                        (mm_interconnect_0_uart_rs_s1_chipselect)                    //                                       .chipselect
	);

	parallel_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_0_irq_irq)                   //    sender.irq
	);

	parallel_irq_mapper_001 irq_mapper_001 (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu_1_irq_irq)                   //    sender.irq
	);

	parallel_irq_mapper_001 irq_mapper_002 (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu_2_irq_irq)                   //    sender.irq
	);

	parallel_irq_mapper_001 irq_mapper_003 (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu_3_irq_irq)                   //    sender.irq
	);

	parallel_irq_mapper_004 irq_mapper_004 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_004_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_receiver0_irq),       // receiver1.irq
		.sender_irq    (hypervisor_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (hypervisor_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_in1      (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

endmodule
